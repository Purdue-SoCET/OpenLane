magic
tech sky130A
magscale 1 2
timestamp 1701386622
<< viali >>
rect 5273 7837 5307 7871
rect 1501 7769 1535 7803
rect 1685 7769 1719 7803
rect 5457 7701 5491 7735
rect 1685 7429 1719 7463
rect 3433 7429 3467 7463
rect 6929 7361 6963 7395
rect 1409 7293 1443 7327
rect 3157 7157 3191 7191
rect 4905 7157 4939 7191
rect 6837 7157 6871 7191
rect 4740 6817 4774 6851
rect 7021 6817 7055 6851
rect 3157 6749 3191 6783
rect 4077 6749 4111 6783
rect 4169 6749 4203 6783
rect 4261 6749 4295 6783
rect 4445 6749 4479 6783
rect 4537 6749 4571 6783
rect 4997 6749 5031 6783
rect 4813 6681 4847 6715
rect 5273 6681 5307 6715
rect 1869 6613 1903 6647
rect 3801 6613 3835 6647
rect 4629 6613 4663 6647
rect 2605 6409 2639 6443
rect 4813 6409 4847 6443
rect 5733 6409 5767 6443
rect 3341 6341 3375 6375
rect 5149 6341 5183 6375
rect 5365 6341 5399 6375
rect 1409 6273 1443 6307
rect 1777 6273 1811 6307
rect 2145 6273 2179 6307
rect 2421 6273 2455 6307
rect 2513 6273 2547 6307
rect 2789 6273 2823 6307
rect 2973 6273 3007 6307
rect 5457 6273 5491 6307
rect 5917 6273 5951 6307
rect 3065 6205 3099 6239
rect 4997 6137 5031 6171
rect 1961 6069 1995 6103
rect 2237 6069 2271 6103
rect 5181 6069 5215 6103
rect 5549 6069 5583 6103
rect 3249 5865 3283 5899
rect 3433 5865 3467 5899
rect 3801 5865 3835 5899
rect 3985 5865 4019 5899
rect 4813 5865 4847 5899
rect 6561 5865 6595 5899
rect 4261 5797 4295 5831
rect 5181 5797 5215 5831
rect 1409 5729 1443 5763
rect 1685 5729 1719 5763
rect 3157 5729 3191 5763
rect 4261 5661 4295 5695
rect 4521 5655 4555 5689
rect 4629 5661 4663 5695
rect 4813 5661 4847 5695
rect 4905 5661 4939 5695
rect 5273 5661 5307 5695
rect 3401 5593 3435 5627
rect 3617 5593 3651 5627
rect 4169 5593 4203 5627
rect 5181 5593 5215 5627
rect 3969 5525 4003 5559
rect 4445 5525 4479 5559
rect 4997 5525 5031 5559
rect 4721 5321 4755 5355
rect 1961 5253 1995 5287
rect 5273 5253 5307 5287
rect 6545 5253 6579 5287
rect 6745 5253 6779 5287
rect 4353 5185 4387 5219
rect 4537 5185 4571 5219
rect 4905 5185 4939 5219
rect 5089 5185 5123 5219
rect 4813 5117 4847 5151
rect 5917 5117 5951 5151
rect 6193 5117 6227 5151
rect 6377 5049 6411 5083
rect 1685 4981 1719 5015
rect 6561 4981 6595 5015
rect 1501 4777 1535 4811
rect 7021 4777 7055 4811
rect 2697 4709 2731 4743
rect 3525 4709 3559 4743
rect 2237 4641 2271 4675
rect 3249 4641 3283 4675
rect 4629 4641 4663 4675
rect 4813 4641 4847 4675
rect 5273 4641 5307 4675
rect 5549 4641 5583 4675
rect 1777 4573 1811 4607
rect 2329 4573 2363 4607
rect 3157 4573 3191 4607
rect 4997 4573 5031 4607
rect 5089 4573 5123 4607
rect 4537 4505 4571 4539
rect 4721 4437 4755 4471
rect 2237 4233 2271 4267
rect 5365 4233 5399 4267
rect 4077 4165 4111 4199
rect 4997 4165 5031 4199
rect 1409 4097 1443 4131
rect 1869 4097 1903 4131
rect 2513 4097 2547 4131
rect 3157 4097 3191 4131
rect 3801 4097 3835 4131
rect 3893 4097 3927 4131
rect 4261 4097 4295 4131
rect 4537 4097 4571 4131
rect 4629 4097 4663 4131
rect 5273 4097 5307 4131
rect 6377 4097 6411 4131
rect 6561 4097 6595 4131
rect 1961 4029 1995 4063
rect 2605 4029 2639 4063
rect 5733 4029 5767 4063
rect 5825 4029 5859 4063
rect 6009 4029 6043 4063
rect 6745 4029 6779 4063
rect 1593 3961 1627 3995
rect 2881 3961 2915 3995
rect 4629 3961 4663 3995
rect 5089 3961 5123 3995
rect 2421 3893 2455 3927
rect 3065 3893 3099 3927
rect 3249 3893 3283 3927
rect 4077 3893 4111 3927
rect 2697 3689 2731 3723
rect 3893 3689 3927 3723
rect 4169 3689 4203 3723
rect 4905 3689 4939 3723
rect 5549 3689 5583 3723
rect 6009 3689 6043 3723
rect 1593 3621 1627 3655
rect 2513 3621 2547 3655
rect 4629 3621 4663 3655
rect 1869 3553 1903 3587
rect 1961 3553 1995 3587
rect 2329 3553 2363 3587
rect 2697 3553 2731 3587
rect 3617 3553 3651 3587
rect 5089 3553 5123 3587
rect 5733 3553 5767 3587
rect 7021 3553 7055 3587
rect 1409 3485 1443 3519
rect 2237 3485 2271 3519
rect 2605 3485 2639 3519
rect 3065 3485 3099 3519
rect 3157 3485 3191 3519
rect 3341 3485 3375 3519
rect 3433 3485 3467 3519
rect 3801 3485 3835 3519
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 4353 3485 4387 3519
rect 4997 3485 5031 3519
rect 5181 3485 5215 3519
rect 5457 3485 5491 3519
rect 6745 3485 6779 3519
rect 4721 3417 4755 3451
rect 2973 3349 3007 3383
rect 5273 3349 5307 3383
rect 2697 3145 2731 3179
rect 3801 3145 3835 3179
rect 4445 3145 4479 3179
rect 5089 3145 5123 3179
rect 5733 3145 5767 3179
rect 6101 3145 6135 3179
rect 1409 3009 1443 3043
rect 2237 3009 2271 3043
rect 2973 3009 3007 3043
rect 3985 3009 4019 3043
rect 4169 3009 4203 3043
rect 4261 3009 4295 3043
rect 4629 3009 4663 3043
rect 4721 3009 4755 3043
rect 4813 3009 4847 3043
rect 4905 3009 4939 3043
rect 5089 3009 5123 3043
rect 5273 3009 5307 3043
rect 5825 3009 5859 3043
rect 5917 3009 5951 3043
rect 6837 3009 6871 3043
rect 3433 2941 3467 2975
rect 6377 2941 6411 2975
rect 2605 2873 2639 2907
rect 1593 2805 1627 2839
rect 3065 2805 3099 2839
rect 6561 2805 6595 2839
rect 6653 2601 6687 2635
rect 6837 2397 6871 2431
rect 6929 2397 6963 2431
rect 6653 2329 6687 2363
<< metal1 >>
rect 1104 8186 7360 8208
rect 1104 8134 2350 8186
rect 2402 8134 2414 8186
rect 2466 8134 2478 8186
rect 2530 8134 2542 8186
rect 2594 8134 2606 8186
rect 2658 8134 7360 8186
rect 1104 8112 7360 8134
rect 5166 7828 5172 7880
rect 5224 7868 5230 7880
rect 5261 7871 5319 7877
rect 5261 7868 5273 7871
rect 5224 7840 5273 7868
rect 5224 7828 5230 7840
rect 5261 7837 5273 7840
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 1486 7760 1492 7812
rect 1544 7760 1550 7812
rect 1673 7803 1731 7809
rect 1673 7769 1685 7803
rect 1719 7800 1731 7803
rect 2130 7800 2136 7812
rect 1719 7772 2136 7800
rect 1719 7769 1731 7772
rect 1673 7763 1731 7769
rect 2130 7760 2136 7772
rect 2188 7800 2194 7812
rect 3878 7800 3884 7812
rect 2188 7772 3884 7800
rect 2188 7760 2194 7772
rect 3878 7760 3884 7772
rect 3936 7760 3942 7812
rect 5442 7692 5448 7744
rect 5500 7692 5506 7744
rect 1104 7642 7360 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 7360 7642
rect 1104 7568 7360 7590
rect 1302 7488 1308 7540
rect 1360 7528 1366 7540
rect 1360 7500 3464 7528
rect 1360 7488 1366 7500
rect 1673 7463 1731 7469
rect 1673 7429 1685 7463
rect 1719 7460 1731 7463
rect 1946 7460 1952 7472
rect 1719 7432 1952 7460
rect 1719 7429 1731 7432
rect 1673 7423 1731 7429
rect 1946 7420 1952 7432
rect 2004 7420 2010 7472
rect 2130 7420 2136 7472
rect 2188 7420 2194 7472
rect 3436 7469 3464 7500
rect 3421 7463 3479 7469
rect 3421 7429 3433 7463
rect 3467 7429 3479 7463
rect 3421 7423 3479 7429
rect 6914 7352 6920 7404
rect 6972 7352 6978 7404
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7293 1455 7327
rect 1397 7287 1455 7293
rect 1412 7188 1440 7287
rect 1854 7188 1860 7200
rect 1412 7160 1860 7188
rect 1854 7148 1860 7160
rect 1912 7148 1918 7200
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 3145 7191 3203 7197
rect 3145 7188 3157 7191
rect 2832 7160 3157 7188
rect 2832 7148 2838 7160
rect 3145 7157 3157 7160
rect 3191 7157 3203 7191
rect 3145 7151 3203 7157
rect 4893 7191 4951 7197
rect 4893 7157 4905 7191
rect 4939 7188 4951 7191
rect 5258 7188 5264 7200
rect 4939 7160 5264 7188
rect 4939 7157 4951 7160
rect 4893 7151 4951 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 6822 7148 6828 7200
rect 6880 7148 6886 7200
rect 1104 7098 7360 7120
rect 1104 7046 2350 7098
rect 2402 7046 2414 7098
rect 2466 7046 2478 7098
rect 2530 7046 2542 7098
rect 2594 7046 2606 7098
rect 2658 7046 7360 7098
rect 1104 7024 7360 7046
rect 2498 6944 2504 6996
rect 2556 6984 2562 6996
rect 4154 6984 4160 6996
rect 2556 6956 4160 6984
rect 2556 6944 2562 6956
rect 4154 6944 4160 6956
rect 4212 6944 4218 6996
rect 4080 6888 4844 6916
rect 4080 6848 4108 6888
rect 4728 6851 4786 6857
rect 4728 6848 4740 6851
rect 3160 6820 4108 6848
rect 4172 6820 4568 6848
rect 3160 6789 3188 6820
rect 4172 6792 4200 6820
rect 4540 6792 4568 6820
rect 4632 6820 4740 6848
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6749 3203 6783
rect 4065 6783 4123 6789
rect 4065 6774 4077 6783
rect 3145 6743 3203 6749
rect 4060 6749 4077 6774
rect 4111 6749 4123 6783
rect 4060 6743 4123 6749
rect 2590 6712 2596 6724
rect 1872 6684 2596 6712
rect 1872 6656 1900 6684
rect 2590 6672 2596 6684
rect 2648 6672 2654 6724
rect 4060 6712 4088 6743
rect 4154 6740 4160 6792
rect 4212 6740 4218 6792
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6777 4307 6783
rect 4295 6749 4384 6777
rect 4249 6743 4307 6749
rect 4356 6712 4384 6749
rect 4430 6740 4436 6792
rect 4488 6740 4494 6792
rect 4522 6740 4528 6792
rect 4580 6740 4586 6792
rect 4632 6712 4660 6820
rect 4728 6817 4740 6820
rect 4774 6817 4786 6851
rect 4816 6848 4844 6888
rect 5258 6848 5264 6860
rect 4816 6820 5264 6848
rect 4728 6811 4786 6817
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 5350 6808 5356 6860
rect 5408 6848 5414 6860
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 5408 6820 7021 6848
rect 5408 6808 5414 6820
rect 7009 6817 7021 6820
rect 7055 6817 7067 6851
rect 7009 6811 7067 6817
rect 4982 6740 4988 6792
rect 5040 6740 5046 6792
rect 4060 6684 4200 6712
rect 4356 6684 4660 6712
rect 4801 6715 4859 6721
rect 1854 6604 1860 6656
rect 1912 6604 1918 6656
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 3476 6616 3801 6644
rect 3476 6604 3482 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 4172 6644 4200 6684
rect 4801 6681 4813 6715
rect 4847 6681 4859 6715
rect 4801 6675 4859 6681
rect 5261 6715 5319 6721
rect 5261 6681 5273 6715
rect 5307 6712 5319 6715
rect 5534 6712 5540 6724
rect 5307 6684 5540 6712
rect 5307 6681 5319 6684
rect 5261 6675 5319 6681
rect 4614 6644 4620 6656
rect 4172 6616 4620 6644
rect 3789 6607 3847 6613
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 4816 6644 4844 6675
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 5994 6672 6000 6724
rect 6052 6672 6058 6724
rect 5442 6644 5448 6656
rect 4816 6616 5448 6644
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 1104 6554 7360 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 7360 6554
rect 1104 6480 7360 6502
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 2593 6443 2651 6449
rect 2593 6440 2605 6443
rect 2188 6412 2605 6440
rect 2188 6400 2194 6412
rect 2593 6409 2605 6412
rect 2639 6440 2651 6443
rect 4614 6440 4620 6452
rect 2639 6412 4620 6440
rect 2639 6409 2651 6412
rect 2593 6403 2651 6409
rect 4614 6400 4620 6412
rect 4672 6440 4678 6452
rect 4801 6443 4859 6449
rect 4801 6440 4813 6443
rect 4672 6412 4813 6440
rect 4672 6400 4678 6412
rect 4801 6409 4813 6412
rect 4847 6409 4859 6443
rect 4801 6403 4859 6409
rect 4890 6400 4896 6452
rect 4948 6440 4954 6452
rect 4948 6412 5396 6440
rect 4948 6400 4954 6412
rect 5368 6384 5396 6412
rect 5442 6400 5448 6452
rect 5500 6400 5506 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 5721 6443 5779 6449
rect 5721 6440 5733 6443
rect 5592 6412 5733 6440
rect 5592 6400 5598 6412
rect 5721 6409 5733 6412
rect 5767 6409 5779 6443
rect 5721 6403 5779 6409
rect 3234 6372 3240 6384
rect 2148 6344 3240 6372
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 2148 6313 2176 6344
rect 3234 6332 3240 6344
rect 3292 6332 3298 6384
rect 3329 6375 3387 6381
rect 3329 6341 3341 6375
rect 3375 6372 3387 6375
rect 3418 6372 3424 6384
rect 3375 6344 3424 6372
rect 3375 6341 3387 6344
rect 3329 6335 3387 6341
rect 3418 6332 3424 6344
rect 3476 6332 3482 6384
rect 4706 6332 4712 6384
rect 4764 6372 4770 6384
rect 5137 6375 5195 6381
rect 5137 6372 5149 6375
rect 4764 6344 5149 6372
rect 4764 6332 4770 6344
rect 5137 6341 5149 6344
rect 5183 6341 5195 6375
rect 5137 6335 5195 6341
rect 5350 6332 5356 6384
rect 5408 6332 5414 6384
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 992 6276 1409 6304
rect 992 6264 998 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 2409 6307 2467 6313
rect 2409 6273 2421 6307
rect 2455 6273 2467 6307
rect 2409 6267 2467 6273
rect 1780 6168 1808 6267
rect 2424 6168 2452 6267
rect 2498 6264 2504 6316
rect 2556 6264 2562 6316
rect 2774 6264 2780 6316
rect 2832 6264 2838 6316
rect 2958 6264 2964 6316
rect 3016 6264 3022 6316
rect 5460 6313 5488 6400
rect 5445 6307 5503 6313
rect 4462 6290 5120 6304
rect 4448 6276 5120 6290
rect 2590 6196 2596 6248
rect 2648 6236 2654 6248
rect 3053 6239 3111 6245
rect 3053 6236 3065 6239
rect 2648 6208 3065 6236
rect 2648 6196 2654 6208
rect 3053 6205 3065 6208
rect 3099 6205 3111 6239
rect 3053 6199 3111 6205
rect 3878 6196 3884 6248
rect 3936 6236 3942 6248
rect 4448 6236 4476 6276
rect 3936 6208 4476 6236
rect 3936 6196 3942 6208
rect 4522 6196 4528 6248
rect 4580 6236 4586 6248
rect 4580 6208 5028 6236
rect 4580 6196 4586 6208
rect 5000 6177 5028 6208
rect 4985 6171 5043 6177
rect 1780 6140 2360 6168
rect 2424 6140 3188 6168
rect 1946 6060 1952 6112
rect 2004 6060 2010 6112
rect 2222 6060 2228 6112
rect 2280 6060 2286 6112
rect 2332 6100 2360 6140
rect 3050 6100 3056 6112
rect 2332 6072 3056 6100
rect 3050 6060 3056 6072
rect 3108 6060 3114 6112
rect 3160 6100 3188 6140
rect 4985 6137 4997 6171
rect 5031 6137 5043 6171
rect 5092 6168 5120 6276
rect 5445 6273 5457 6307
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5902 6264 5908 6316
rect 5960 6264 5966 6316
rect 5994 6168 6000 6180
rect 5092 6140 6000 6168
rect 4985 6131 5043 6137
rect 5994 6128 6000 6140
rect 6052 6128 6058 6180
rect 3786 6100 3792 6112
rect 3160 6072 3792 6100
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 5169 6103 5227 6109
rect 5169 6100 5181 6103
rect 4028 6072 5181 6100
rect 4028 6060 4034 6072
rect 5169 6069 5181 6072
rect 5215 6069 5227 6103
rect 5169 6063 5227 6069
rect 5350 6060 5356 6112
rect 5408 6100 5414 6112
rect 5537 6103 5595 6109
rect 5537 6100 5549 6103
rect 5408 6072 5549 6100
rect 5408 6060 5414 6072
rect 5537 6069 5549 6072
rect 5583 6069 5595 6103
rect 5537 6063 5595 6069
rect 1104 6010 7360 6032
rect 1104 5958 2350 6010
rect 2402 5958 2414 6010
rect 2466 5958 2478 6010
rect 2530 5958 2542 6010
rect 2594 5958 2606 6010
rect 2658 5958 7360 6010
rect 1104 5936 7360 5958
rect 1854 5896 1860 5908
rect 1412 5868 1860 5896
rect 1412 5769 1440 5868
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 3234 5856 3240 5908
rect 3292 5856 3298 5908
rect 3421 5899 3479 5905
rect 3421 5865 3433 5899
rect 3467 5865 3479 5899
rect 3421 5859 3479 5865
rect 3436 5828 3464 5859
rect 3786 5856 3792 5908
rect 3844 5856 3850 5908
rect 3973 5899 4031 5905
rect 3973 5865 3985 5899
rect 4019 5896 4031 5899
rect 4430 5896 4436 5908
rect 4019 5868 4436 5896
rect 4019 5865 4031 5868
rect 3973 5859 4031 5865
rect 3988 5828 4016 5859
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 4522 5856 4528 5908
rect 4580 5856 4586 5908
rect 4614 5856 4620 5908
rect 4672 5896 4678 5908
rect 4801 5899 4859 5905
rect 4801 5896 4813 5899
rect 4672 5868 4813 5896
rect 4672 5856 4678 5868
rect 4801 5865 4813 5868
rect 4847 5865 4859 5899
rect 6549 5899 6607 5905
rect 6549 5896 6561 5899
rect 4801 5859 4859 5865
rect 5000 5868 6561 5896
rect 3436 5800 4016 5828
rect 4249 5831 4307 5837
rect 4249 5797 4261 5831
rect 4295 5797 4307 5831
rect 4540 5828 4568 5856
rect 5000 5840 5028 5868
rect 6549 5865 6561 5868
rect 6595 5865 6607 5899
rect 6549 5859 6607 5865
rect 4540 5800 4844 5828
rect 4249 5791 4307 5797
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5729 1455 5763
rect 1397 5723 1455 5729
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5760 1731 5763
rect 2222 5760 2228 5772
rect 1719 5732 2228 5760
rect 1719 5729 1731 5732
rect 1673 5723 1731 5729
rect 2222 5720 2228 5732
rect 2280 5720 2286 5772
rect 3050 5720 3056 5772
rect 3108 5760 3114 5772
rect 3145 5763 3203 5769
rect 3145 5760 3157 5763
rect 3108 5732 3157 5760
rect 3108 5720 3114 5732
rect 3145 5729 3157 5732
rect 3191 5760 3203 5763
rect 3510 5760 3516 5772
rect 3191 5732 3516 5760
rect 3191 5729 3203 5732
rect 3145 5723 3203 5729
rect 3510 5720 3516 5732
rect 3568 5760 3574 5772
rect 3970 5760 3976 5772
rect 3568 5732 3976 5760
rect 3568 5720 3574 5732
rect 3970 5720 3976 5732
rect 4028 5760 4034 5772
rect 4264 5760 4292 5791
rect 4028 5732 4200 5760
rect 4264 5732 4771 5760
rect 4028 5720 4034 5732
rect 3878 5692 3884 5704
rect 2806 5664 3884 5692
rect 3878 5652 3884 5664
rect 3936 5652 3942 5704
rect 4172 5692 4200 5732
rect 4249 5695 4307 5701
rect 4249 5692 4261 5695
rect 4172 5664 4261 5692
rect 4249 5661 4261 5664
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 4338 5652 4344 5704
rect 4396 5692 4402 5704
rect 4617 5695 4675 5701
rect 4396 5686 4476 5692
rect 4509 5689 4567 5695
rect 4509 5686 4521 5689
rect 4396 5664 4521 5686
rect 4396 5652 4402 5664
rect 4448 5658 4521 5664
rect 4509 5655 4521 5658
rect 4555 5655 4567 5689
rect 4617 5661 4629 5695
rect 4663 5686 4675 5695
rect 4743 5686 4771 5732
rect 4816 5701 4844 5800
rect 4982 5788 4988 5840
rect 5040 5788 5046 5840
rect 5169 5831 5227 5837
rect 5169 5797 5181 5831
rect 5215 5828 5227 5831
rect 5534 5828 5540 5840
rect 5215 5800 5540 5828
rect 5215 5797 5227 5800
rect 5169 5791 5227 5797
rect 5534 5788 5540 5800
rect 5592 5788 5598 5840
rect 4663 5661 4771 5686
rect 4617 5658 4771 5661
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5661 4859 5695
rect 4617 5655 4675 5658
rect 4801 5655 4859 5661
rect 4509 5649 4567 5655
rect 4890 5652 4896 5704
rect 4948 5652 4954 5704
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 5442 5652 5448 5704
rect 5500 5652 5506 5704
rect 2958 5584 2964 5636
rect 3016 5624 3022 5636
rect 3389 5627 3447 5633
rect 3389 5624 3401 5627
rect 3016 5596 3401 5624
rect 3016 5584 3022 5596
rect 3389 5593 3401 5596
rect 3435 5593 3447 5627
rect 3389 5587 3447 5593
rect 3605 5627 3663 5633
rect 3605 5593 3617 5627
rect 3651 5624 3663 5627
rect 4154 5624 4160 5636
rect 3651 5596 4160 5624
rect 3651 5593 3663 5596
rect 3605 5587 3663 5593
rect 4154 5584 4160 5596
rect 4212 5584 4218 5636
rect 5169 5627 5227 5633
rect 5169 5593 5181 5627
rect 5215 5624 5227 5627
rect 5460 5624 5488 5652
rect 5215 5596 5488 5624
rect 5215 5593 5227 5596
rect 5169 5587 5227 5593
rect 3957 5559 4015 5565
rect 3957 5525 3969 5559
rect 4003 5556 4015 5559
rect 4062 5556 4068 5568
rect 4003 5528 4068 5556
rect 4003 5525 4015 5528
rect 3957 5519 4015 5525
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 4433 5559 4491 5565
rect 4433 5525 4445 5559
rect 4479 5556 4491 5559
rect 4706 5556 4712 5568
rect 4479 5528 4712 5556
rect 4479 5525 4491 5528
rect 4433 5519 4491 5525
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 4985 5559 5043 5565
rect 4985 5556 4997 5559
rect 4856 5528 4997 5556
rect 4856 5516 4862 5528
rect 4985 5525 4997 5528
rect 5031 5525 5043 5559
rect 4985 5519 5043 5525
rect 1104 5466 7360 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 7360 5466
rect 1104 5392 7360 5414
rect 4338 5312 4344 5364
rect 4396 5352 4402 5364
rect 4614 5352 4620 5364
rect 4396 5324 4620 5352
rect 4396 5312 4402 5324
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 4709 5355 4767 5361
rect 4709 5321 4721 5355
rect 4755 5352 4767 5355
rect 4798 5352 4804 5364
rect 4755 5324 4804 5352
rect 4755 5321 4767 5324
rect 4709 5315 4767 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5074 5312 5080 5364
rect 5132 5352 5138 5364
rect 5132 5324 6776 5352
rect 5132 5312 5138 5324
rect 1949 5287 2007 5293
rect 1949 5253 1961 5287
rect 1995 5284 2007 5287
rect 2866 5284 2872 5296
rect 1995 5256 2872 5284
rect 1995 5253 2007 5256
rect 1949 5247 2007 5253
rect 2866 5244 2872 5256
rect 2924 5244 2930 5296
rect 4154 5244 4160 5296
rect 4212 5284 4218 5296
rect 6748 5293 6776 5324
rect 5261 5287 5319 5293
rect 4212 5256 5120 5284
rect 4212 5244 4218 5256
rect 4338 5176 4344 5228
rect 4396 5176 4402 5228
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 4540 5080 4568 5179
rect 4614 5176 4620 5228
rect 4672 5216 4678 5228
rect 5092 5225 5120 5256
rect 5261 5253 5273 5287
rect 5307 5284 5319 5287
rect 6533 5287 6591 5293
rect 6533 5284 6545 5287
rect 5307 5256 6545 5284
rect 5307 5253 5319 5256
rect 5261 5247 5319 5253
rect 6533 5253 6545 5256
rect 6579 5284 6591 5287
rect 6733 5287 6791 5293
rect 6579 5256 6684 5284
rect 6579 5253 6591 5256
rect 6533 5247 6591 5253
rect 6656 5228 6684 5256
rect 6733 5253 6745 5287
rect 6779 5253 6791 5287
rect 6733 5247 6791 5253
rect 4893 5219 4951 5225
rect 4893 5216 4905 5219
rect 4672 5188 4905 5216
rect 4672 5176 4678 5188
rect 4893 5185 4905 5188
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 5350 5216 5356 5228
rect 5123 5188 5356 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 4706 5108 4712 5160
rect 4764 5148 4770 5160
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 4764 5120 4813 5148
rect 4764 5108 4770 5120
rect 4801 5117 4813 5120
rect 4847 5117 4859 5151
rect 4908 5148 4936 5179
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 6638 5176 6644 5228
rect 6696 5176 6702 5228
rect 5258 5148 5264 5160
rect 4908 5120 5264 5148
rect 4801 5111 4859 5117
rect 5258 5108 5264 5120
rect 5316 5148 5322 5160
rect 5905 5151 5963 5157
rect 5905 5148 5917 5151
rect 5316 5120 5917 5148
rect 5316 5108 5322 5120
rect 5905 5117 5917 5120
rect 5951 5117 5963 5151
rect 5905 5111 5963 5117
rect 6181 5151 6239 5157
rect 6181 5117 6193 5151
rect 6227 5148 6239 5151
rect 7006 5148 7012 5160
rect 6227 5120 7012 5148
rect 6227 5117 6239 5120
rect 6181 5111 6239 5117
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 5074 5080 5080 5092
rect 4540 5052 5080 5080
rect 5074 5040 5080 5052
rect 5132 5040 5138 5092
rect 5166 5040 5172 5092
rect 5224 5080 5230 5092
rect 6365 5083 6423 5089
rect 6365 5080 6377 5083
rect 5224 5052 6377 5080
rect 5224 5040 5230 5052
rect 6365 5049 6377 5052
rect 6411 5049 6423 5083
rect 6365 5043 6423 5049
rect 934 4972 940 5024
rect 992 5012 998 5024
rect 1673 5015 1731 5021
rect 1673 5012 1685 5015
rect 992 4984 1685 5012
rect 992 4972 998 4984
rect 1673 4981 1685 4984
rect 1719 4981 1731 5015
rect 1673 4975 1731 4981
rect 6549 5015 6607 5021
rect 6549 4981 6561 5015
rect 6595 5012 6607 5015
rect 6822 5012 6828 5024
rect 6595 4984 6828 5012
rect 6595 4981 6607 4984
rect 6549 4975 6607 4981
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 1104 4922 7360 4944
rect 1104 4870 2350 4922
rect 2402 4870 2414 4922
rect 2466 4870 2478 4922
rect 2530 4870 2542 4922
rect 2594 4870 2606 4922
rect 2658 4870 7360 4922
rect 1104 4848 7360 4870
rect 1026 4768 1032 4820
rect 1084 4808 1090 4820
rect 1489 4811 1547 4817
rect 1489 4808 1501 4811
rect 1084 4780 1501 4808
rect 1084 4768 1090 4780
rect 1489 4777 1501 4780
rect 1535 4777 1547 4811
rect 1489 4771 1547 4777
rect 4982 4768 4988 4820
rect 5040 4768 5046 4820
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7009 4811 7067 4817
rect 7009 4808 7021 4811
rect 6972 4780 7021 4808
rect 6972 4768 6978 4780
rect 7009 4777 7021 4780
rect 7055 4777 7067 4811
rect 7009 4771 7067 4777
rect 2685 4743 2743 4749
rect 2685 4709 2697 4743
rect 2731 4740 2743 4743
rect 3513 4743 3571 4749
rect 2731 4712 3464 4740
rect 2731 4709 2743 4712
rect 2685 4703 2743 4709
rect 2222 4632 2228 4684
rect 2280 4632 2286 4684
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4672 3295 4675
rect 3326 4672 3332 4684
rect 3283 4644 3332 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 3436 4672 3464 4712
rect 3513 4709 3525 4743
rect 3559 4740 3571 4743
rect 3559 4712 4844 4740
rect 3559 4709 3571 4712
rect 3513 4703 3571 4709
rect 4816 4681 4844 4712
rect 4617 4675 4675 4681
rect 4617 4672 4629 4675
rect 3436 4644 4629 4672
rect 4617 4641 4629 4644
rect 4663 4641 4675 4675
rect 4617 4635 4675 4641
rect 4801 4675 4859 4681
rect 4801 4641 4813 4675
rect 4847 4641 4859 4675
rect 5000 4672 5028 4768
rect 5261 4675 5319 4681
rect 5261 4672 5273 4675
rect 5000 4644 5273 4672
rect 4801 4635 4859 4641
rect 5261 4641 5273 4644
rect 5307 4641 5319 4675
rect 5261 4635 5319 4641
rect 5534 4632 5540 4684
rect 5592 4632 5598 4684
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 2130 4604 2136 4616
rect 1811 4576 2136 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 2314 4564 2320 4616
rect 2372 4564 2378 4616
rect 2774 4564 2780 4616
rect 2832 4604 2838 4616
rect 3145 4607 3203 4613
rect 3145 4604 3157 4607
rect 2832 4576 3157 4604
rect 2832 4564 2838 4576
rect 3145 4573 3157 4576
rect 3191 4573 3203 4607
rect 3145 4567 3203 4573
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4573 5043 4607
rect 4985 4567 5043 4573
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4604 5135 4607
rect 5166 4604 5172 4616
rect 5123 4576 5172 4604
rect 5123 4573 5135 4576
rect 5077 4567 5135 4573
rect 2148 4536 2176 4564
rect 3602 4536 3608 4548
rect 2148 4508 3608 4536
rect 3602 4496 3608 4508
rect 3660 4496 3666 4548
rect 4525 4539 4583 4545
rect 4525 4505 4537 4539
rect 4571 4536 4583 4539
rect 4890 4536 4896 4548
rect 4571 4508 4896 4536
rect 4571 4505 4583 4508
rect 4525 4499 4583 4505
rect 4890 4496 4896 4508
rect 4948 4496 4954 4548
rect 5000 4536 5028 4567
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 5810 4536 5816 4548
rect 5000 4508 5816 4536
rect 5810 4496 5816 4508
rect 5868 4496 5874 4548
rect 5994 4496 6000 4548
rect 6052 4496 6058 4548
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4709 4471 4767 4477
rect 4709 4468 4721 4471
rect 4212 4440 4721 4468
rect 4212 4428 4218 4440
rect 4709 4437 4721 4440
rect 4755 4437 4767 4471
rect 4709 4431 4767 4437
rect 1104 4378 7360 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 7360 4378
rect 1104 4304 7360 4326
rect 2225 4267 2283 4273
rect 2225 4233 2237 4267
rect 2271 4264 2283 4267
rect 4154 4264 4160 4276
rect 2271 4236 4160 4264
rect 2271 4233 2283 4236
rect 2225 4227 2283 4233
rect 4154 4224 4160 4236
rect 4212 4224 4218 4276
rect 5258 4224 5264 4276
rect 5316 4264 5322 4276
rect 5353 4267 5411 4273
rect 5353 4264 5365 4267
rect 5316 4236 5365 4264
rect 5316 4224 5322 4236
rect 5353 4233 5365 4236
rect 5399 4233 5411 4267
rect 5353 4227 5411 4233
rect 2682 4196 2688 4208
rect 2516 4168 2688 4196
rect 1394 4088 1400 4140
rect 1452 4088 1458 4140
rect 1854 4088 1860 4140
rect 1912 4088 1918 4140
rect 2516 4137 2544 4168
rect 2682 4156 2688 4168
rect 2740 4156 2746 4208
rect 4065 4199 4123 4205
rect 4065 4165 4077 4199
rect 4111 4165 4123 4199
rect 4985 4199 5043 4205
rect 4065 4159 4123 4165
rect 4540 4168 4752 4196
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4097 2559 4131
rect 2501 4091 2559 4097
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 3145 4131 3203 4137
rect 3145 4128 3157 4131
rect 2832 4100 3157 4128
rect 2832 4088 2838 4100
rect 3145 4097 3157 4100
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3786 4088 3792 4140
rect 3844 4088 3850 4140
rect 3878 4088 3884 4140
rect 3936 4088 3942 4140
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4080 4128 4108 4159
rect 4028 4100 4108 4128
rect 4028 4088 4034 4100
rect 4246 4088 4252 4140
rect 4304 4088 4310 4140
rect 4540 4137 4568 4168
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4724 4128 4752 4168
rect 4985 4165 4997 4199
rect 5031 4196 5043 4199
rect 5276 4196 5304 4224
rect 5031 4168 5304 4196
rect 5031 4165 5043 4168
rect 4985 4159 5043 4165
rect 5261 4131 5319 4137
rect 4724 4100 4844 4128
rect 4617 4091 4675 4097
rect 1946 4020 1952 4072
rect 2004 4020 2010 4072
rect 2593 4063 2651 4069
rect 2593 4029 2605 4063
rect 2639 4060 2651 4063
rect 3510 4060 3516 4072
rect 2639 4032 3516 4060
rect 2639 4029 2651 4032
rect 2593 4023 2651 4029
rect 3510 4020 3516 4032
rect 3568 4020 3574 4072
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 4632 4060 4660 4091
rect 4120 4032 4660 4060
rect 4816 4060 4844 4100
rect 5261 4097 5273 4131
rect 5307 4128 5319 4131
rect 5307 4100 5488 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 4816 4032 5120 4060
rect 4120 4020 4126 4032
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 2774 3992 2780 4004
rect 1627 3964 2780 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 2774 3952 2780 3964
rect 2832 3952 2838 4004
rect 2869 3995 2927 4001
rect 2869 3961 2881 3995
rect 2915 3961 2927 3995
rect 4338 3992 4344 4004
rect 2869 3955 2927 3961
rect 2976 3964 4344 3992
rect 2222 3884 2228 3936
rect 2280 3924 2286 3936
rect 2409 3927 2467 3933
rect 2409 3924 2421 3927
rect 2280 3896 2421 3924
rect 2280 3884 2286 3896
rect 2409 3893 2421 3896
rect 2455 3893 2467 3927
rect 2409 3887 2467 3893
rect 2498 3884 2504 3936
rect 2556 3924 2562 3936
rect 2884 3924 2912 3955
rect 2976 3936 3004 3964
rect 4338 3952 4344 3964
rect 4396 3992 4402 4004
rect 4396 3964 4568 3992
rect 4396 3952 4402 3964
rect 2556 3896 2912 3924
rect 2556 3884 2562 3896
rect 2958 3884 2964 3936
rect 3016 3884 3022 3936
rect 3050 3884 3056 3936
rect 3108 3884 3114 3936
rect 3234 3884 3240 3936
rect 3292 3884 3298 3936
rect 4062 3884 4068 3936
rect 4120 3884 4126 3936
rect 4540 3924 4568 3964
rect 4614 3952 4620 4004
rect 4672 3952 4678 4004
rect 5092 4001 5120 4032
rect 5077 3995 5135 4001
rect 5077 3961 5089 3995
rect 5123 3961 5135 3995
rect 5077 3955 5135 3961
rect 5460 3936 5488 4100
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 5960 4100 6377 4128
rect 5960 4088 5966 4100
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 6638 4128 6644 4140
rect 6595 4100 6644 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 5718 4020 5724 4072
rect 5776 4020 5782 4072
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4029 5871 4063
rect 5813 4023 5871 4029
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4060 6055 4063
rect 6733 4063 6791 4069
rect 6733 4060 6745 4063
rect 6043 4032 6745 4060
rect 6043 4029 6055 4032
rect 5997 4023 6055 4029
rect 6733 4029 6745 4032
rect 6779 4060 6791 4063
rect 6822 4060 6828 4072
rect 6779 4032 6828 4060
rect 6779 4029 6791 4032
rect 6733 4023 6791 4029
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 5828 3992 5856 4023
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 5684 3964 5856 3992
rect 5684 3952 5690 3964
rect 5258 3924 5264 3936
rect 4540 3896 5264 3924
rect 5258 3884 5264 3896
rect 5316 3884 5322 3936
rect 5442 3884 5448 3936
rect 5500 3884 5506 3936
rect 1104 3834 7360 3856
rect 1104 3782 2350 3834
rect 2402 3782 2414 3834
rect 2466 3782 2478 3834
rect 2530 3782 2542 3834
rect 2594 3782 2606 3834
rect 2658 3782 7360 3834
rect 1104 3760 7360 3782
rect 1854 3680 1860 3732
rect 1912 3680 1918 3732
rect 2222 3680 2228 3732
rect 2280 3680 2286 3732
rect 2685 3723 2743 3729
rect 2685 3689 2697 3723
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 1581 3655 1639 3661
rect 1581 3621 1593 3655
rect 1627 3652 1639 3655
rect 1872 3652 1900 3680
rect 1627 3624 1900 3652
rect 1627 3621 1639 3624
rect 1581 3615 1639 3621
rect 1872 3593 1900 3624
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 2240 3584 2268 3680
rect 2501 3655 2559 3661
rect 2501 3621 2513 3655
rect 2547 3652 2559 3655
rect 2590 3652 2596 3664
rect 2547 3624 2596 3652
rect 2547 3621 2559 3624
rect 2501 3615 2559 3621
rect 2590 3612 2596 3624
rect 2648 3612 2654 3664
rect 2700 3652 2728 3683
rect 3878 3680 3884 3732
rect 3936 3680 3942 3732
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 4157 3723 4215 3729
rect 4157 3720 4169 3723
rect 4120 3692 4169 3720
rect 4120 3680 4126 3692
rect 4157 3689 4169 3692
rect 4203 3689 4215 3723
rect 4798 3720 4804 3732
rect 4157 3683 4215 3689
rect 4264 3692 4804 3720
rect 2774 3652 2780 3664
rect 2700 3624 2780 3652
rect 2774 3612 2780 3624
rect 2832 3612 2838 3664
rect 3050 3612 3056 3664
rect 3108 3612 3114 3664
rect 3234 3612 3240 3664
rect 3292 3612 3298 3664
rect 3970 3612 3976 3664
rect 4028 3652 4034 3664
rect 4264 3652 4292 3692
rect 4798 3680 4804 3692
rect 4856 3720 4862 3732
rect 4893 3723 4951 3729
rect 4893 3720 4905 3723
rect 4856 3692 4905 3720
rect 4856 3680 4862 3692
rect 4893 3689 4905 3692
rect 4939 3689 4951 3723
rect 4893 3683 4951 3689
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5534 3720 5540 3732
rect 5132 3692 5540 3720
rect 5132 3680 5138 3692
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 5626 3680 5632 3732
rect 5684 3680 5690 3732
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 5997 3723 6055 3729
rect 5997 3720 6009 3723
rect 5776 3692 6009 3720
rect 5776 3680 5782 3692
rect 5997 3689 6009 3692
rect 6043 3689 6055 3723
rect 5997 3683 6055 3689
rect 4028 3624 4292 3652
rect 4617 3655 4675 3661
rect 4028 3612 4034 3624
rect 4617 3621 4629 3655
rect 4663 3652 4675 3655
rect 5644 3652 5672 3680
rect 4663 3624 5672 3652
rect 4663 3621 4675 3624
rect 4617 3615 4675 3621
rect 1995 3556 2268 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 992 3488 1409 3516
rect 992 3476 998 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 1872 3448 1900 3547
rect 2314 3544 2320 3596
rect 2372 3544 2378 3596
rect 2685 3587 2743 3593
rect 2685 3584 2697 3587
rect 2424 3556 2697 3584
rect 2038 3476 2044 3528
rect 2096 3516 2102 3528
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 2096 3488 2237 3516
rect 2096 3476 2102 3488
rect 2225 3485 2237 3488
rect 2271 3485 2283 3519
rect 2424 3516 2452 3556
rect 2685 3553 2697 3556
rect 2731 3553 2743 3587
rect 3068 3584 3096 3612
rect 3252 3584 3280 3612
rect 3605 3587 3663 3593
rect 3068 3556 3180 3584
rect 3252 3556 3464 3584
rect 2685 3547 2743 3553
rect 2225 3479 2283 3485
rect 2332 3488 2452 3516
rect 2593 3519 2651 3525
rect 2332 3448 2360 3488
rect 2593 3485 2605 3519
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 1872 3420 2360 3448
rect 2240 3392 2268 3420
rect 2498 3408 2504 3460
rect 2556 3448 2562 3460
rect 2608 3448 2636 3479
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3050 3516 3056 3528
rect 2924 3488 3056 3516
rect 2924 3476 2930 3488
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 3152 3525 3180 3556
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 3234 3516 3240 3528
rect 3191 3488 3240 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 3436 3525 3464 3556
rect 3605 3553 3617 3587
rect 3651 3584 3663 3587
rect 4522 3584 4528 3596
rect 3651 3556 4528 3584
rect 3651 3553 3663 3556
rect 3605 3547 3663 3553
rect 4522 3544 4528 3556
rect 4580 3584 4586 3596
rect 5077 3587 5135 3593
rect 5077 3584 5089 3587
rect 4580 3556 5089 3584
rect 4580 3544 4586 3556
rect 5077 3553 5089 3556
rect 5123 3553 5135 3587
rect 5077 3547 5135 3553
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 5721 3587 5779 3593
rect 5721 3584 5733 3587
rect 5316 3556 5733 3584
rect 5316 3544 5322 3556
rect 5721 3553 5733 3556
rect 5767 3553 5779 3587
rect 5721 3547 5779 3553
rect 7006 3544 7012 3596
rect 7064 3544 7070 3596
rect 3329 3519 3387 3525
rect 3329 3485 3341 3519
rect 3375 3485 3387 3519
rect 3329 3479 3387 3485
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3467 3488 3801 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 2556 3420 2636 3448
rect 3344 3448 3372 3479
rect 3602 3448 3608 3460
rect 3344 3420 3608 3448
rect 2556 3408 2562 3420
rect 3602 3408 3608 3420
rect 3660 3448 3666 3460
rect 3988 3448 4016 3479
rect 4062 3476 4068 3528
rect 4120 3476 4126 3528
rect 4246 3476 4252 3528
rect 4304 3516 4310 3528
rect 4341 3519 4399 3525
rect 4341 3516 4353 3519
rect 4304 3488 4353 3516
rect 4304 3476 4310 3488
rect 4341 3485 4353 3488
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 3660 3420 4016 3448
rect 3660 3408 3666 3420
rect 2222 3340 2228 3392
rect 2280 3340 2286 3392
rect 2958 3340 2964 3392
rect 3016 3340 3022 3392
rect 3050 3340 3056 3392
rect 3108 3380 3114 3392
rect 4356 3380 4384 3479
rect 4982 3476 4988 3528
rect 5040 3476 5046 3528
rect 5166 3476 5172 3528
rect 5224 3476 5230 3528
rect 5442 3476 5448 3528
rect 5500 3476 5506 3528
rect 5534 3476 5540 3528
rect 5592 3516 5598 3528
rect 6546 3516 6552 3528
rect 5592 3488 6552 3516
rect 5592 3476 5598 3488
rect 6546 3476 6552 3488
rect 6604 3516 6610 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6604 3488 6745 3516
rect 6604 3476 6610 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 4709 3451 4767 3457
rect 4709 3417 4721 3451
rect 4755 3448 4767 3451
rect 5460 3448 5488 3476
rect 4755 3420 5488 3448
rect 4755 3417 4767 3420
rect 4709 3411 4767 3417
rect 3108 3352 4384 3380
rect 5261 3383 5319 3389
rect 3108 3340 3114 3352
rect 5261 3349 5273 3383
rect 5307 3380 5319 3383
rect 5552 3380 5580 3476
rect 5307 3352 5580 3380
rect 5307 3349 5319 3352
rect 5261 3343 5319 3349
rect 1104 3290 7360 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 7360 3290
rect 1104 3216 7360 3238
rect 2222 3136 2228 3188
rect 2280 3136 2286 3188
rect 2685 3179 2743 3185
rect 2685 3145 2697 3179
rect 2731 3176 2743 3179
rect 2866 3176 2872 3188
rect 2731 3148 2872 3176
rect 2731 3145 2743 3148
rect 2685 3139 2743 3145
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 3418 3136 3424 3188
rect 3476 3136 3482 3188
rect 3786 3136 3792 3188
rect 3844 3136 3850 3188
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 4433 3179 4491 3185
rect 4433 3176 4445 3179
rect 4120 3148 4445 3176
rect 4120 3136 4126 3148
rect 4433 3145 4445 3148
rect 4479 3145 4491 3179
rect 4433 3139 4491 3145
rect 4522 3136 4528 3188
rect 4580 3136 4586 3188
rect 4982 3176 4988 3188
rect 4816 3148 4988 3176
rect 934 3000 940 3052
rect 992 3040 998 3052
rect 2240 3049 2268 3136
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 992 3012 1409 3040
rect 992 3000 998 3012
rect 1397 3009 1409 3012
rect 1443 3009 1455 3043
rect 1397 3003 1455 3009
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3009 3019 3043
rect 3436 3040 3464 3136
rect 4540 3108 4568 3136
rect 4816 3108 4844 3148
rect 4982 3136 4988 3148
rect 5040 3176 5046 3188
rect 5077 3179 5135 3185
rect 5077 3176 5089 3179
rect 5040 3148 5089 3176
rect 5040 3136 5046 3148
rect 5077 3145 5089 3148
rect 5123 3145 5135 3179
rect 5077 3139 5135 3145
rect 5166 3136 5172 3188
rect 5224 3176 5230 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 5224 3148 5733 3176
rect 5224 3136 5230 3148
rect 5721 3145 5733 3148
rect 5767 3145 5779 3179
rect 5721 3139 5779 3145
rect 6089 3179 6147 3185
rect 6089 3145 6101 3179
rect 6135 3176 6147 3179
rect 6914 3176 6920 3188
rect 6135 3148 6920 3176
rect 6135 3145 6147 3148
rect 6089 3139 6147 3145
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 4172 3080 4384 3108
rect 4540 3080 4660 3108
rect 4172 3049 4200 3080
rect 3973 3043 4031 3049
rect 3973 3040 3985 3043
rect 3436 3012 3985 3040
rect 2961 3003 3019 3009
rect 3973 3009 3985 3012
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 2593 2907 2651 2913
rect 2593 2873 2605 2907
rect 2639 2904 2651 2907
rect 2682 2904 2688 2916
rect 2639 2876 2688 2904
rect 2639 2873 2651 2876
rect 2593 2867 2651 2873
rect 2682 2864 2688 2876
rect 2740 2864 2746 2916
rect 2976 2904 3004 3003
rect 3421 2975 3479 2981
rect 3421 2941 3433 2975
rect 3467 2972 3479 2975
rect 4172 2972 4200 3003
rect 3467 2944 4200 2972
rect 3467 2941 3479 2944
rect 3421 2935 3479 2941
rect 3510 2904 3516 2916
rect 2976 2876 3516 2904
rect 3510 2864 3516 2876
rect 3568 2864 3574 2916
rect 4264 2904 4292 3003
rect 4356 2972 4384 3080
rect 4632 3049 4660 3080
rect 4724 3080 4844 3108
rect 5000 3080 5856 3108
rect 4724 3049 4752 3080
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3009 4767 3043
rect 4709 3003 4767 3009
rect 4798 3000 4804 3052
rect 4856 3000 4862 3052
rect 4890 3000 4896 3052
rect 4948 3040 4954 3052
rect 5000 3040 5028 3080
rect 5828 3049 5856 3080
rect 4948 3012 5028 3040
rect 5077 3043 5135 3049
rect 4948 3000 4954 3012
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 5905 3043 5963 3049
rect 5905 3040 5917 3043
rect 5859 3012 5917 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 5905 3009 5917 3012
rect 5951 3040 5963 3043
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 5951 3012 6837 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 5092 2972 5120 3003
rect 4356 2944 5120 2972
rect 5276 2972 5304 3003
rect 6365 2975 6423 2981
rect 6365 2972 6377 2975
rect 5276 2944 6377 2972
rect 5276 2904 5304 2944
rect 6365 2941 6377 2944
rect 6411 2941 6423 2975
rect 6365 2935 6423 2941
rect 4264 2876 5304 2904
rect 1581 2839 1639 2845
rect 1581 2805 1593 2839
rect 1627 2836 1639 2839
rect 2130 2836 2136 2848
rect 1627 2808 2136 2836
rect 1627 2805 1639 2808
rect 1581 2799 1639 2805
rect 2130 2796 2136 2808
rect 2188 2836 2194 2848
rect 2498 2836 2504 2848
rect 2188 2808 2504 2836
rect 2188 2796 2194 2808
rect 2498 2796 2504 2808
rect 2556 2836 2562 2848
rect 3053 2839 3111 2845
rect 3053 2836 3065 2839
rect 2556 2808 3065 2836
rect 2556 2796 2562 2808
rect 3053 2805 3065 2808
rect 3099 2805 3111 2839
rect 3053 2799 3111 2805
rect 6546 2796 6552 2848
rect 6604 2796 6610 2848
rect 1104 2746 7360 2768
rect 1104 2694 2350 2746
rect 2402 2694 2414 2746
rect 2466 2694 2478 2746
rect 2530 2694 2542 2746
rect 2594 2694 2606 2746
rect 2658 2694 7360 2746
rect 1104 2672 7360 2694
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 5868 2604 6653 2632
rect 5868 2592 5874 2604
rect 6641 2601 6653 2604
rect 6687 2601 6699 2635
rect 6641 2595 6699 2601
rect 6638 2456 6644 2508
rect 6696 2496 6702 2508
rect 6696 2468 6960 2496
rect 6696 2456 6702 2468
rect 6546 2388 6552 2440
rect 6604 2388 6610 2440
rect 6822 2388 6828 2440
rect 6880 2388 6886 2440
rect 6932 2437 6960 2468
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 6564 2360 6592 2388
rect 6641 2363 6699 2369
rect 6641 2360 6653 2363
rect 6564 2332 6653 2360
rect 6641 2329 6653 2332
rect 6687 2329 6699 2363
rect 6641 2323 6699 2329
rect 1104 2202 7360 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 7360 2202
rect 1104 2128 7360 2150
<< via1 >>
rect 2350 8134 2402 8186
rect 2414 8134 2466 8186
rect 2478 8134 2530 8186
rect 2542 8134 2594 8186
rect 2606 8134 2658 8186
rect 5172 7828 5224 7880
rect 1492 7803 1544 7812
rect 1492 7769 1501 7803
rect 1501 7769 1535 7803
rect 1535 7769 1544 7803
rect 1492 7760 1544 7769
rect 2136 7760 2188 7812
rect 3884 7760 3936 7812
rect 5448 7735 5500 7744
rect 5448 7701 5457 7735
rect 5457 7701 5491 7735
rect 5491 7701 5500 7735
rect 5448 7692 5500 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 1308 7488 1360 7540
rect 1952 7420 2004 7472
rect 2136 7420 2188 7472
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 1860 7148 1912 7200
rect 2780 7148 2832 7200
rect 5264 7148 5316 7200
rect 6828 7191 6880 7200
rect 6828 7157 6837 7191
rect 6837 7157 6871 7191
rect 6871 7157 6880 7191
rect 6828 7148 6880 7157
rect 2350 7046 2402 7098
rect 2414 7046 2466 7098
rect 2478 7046 2530 7098
rect 2542 7046 2594 7098
rect 2606 7046 2658 7098
rect 2504 6944 2556 6996
rect 4160 6944 4212 6996
rect 2596 6672 2648 6724
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 5264 6808 5316 6860
rect 5356 6808 5408 6860
rect 4988 6783 5040 6792
rect 4988 6749 4997 6783
rect 4997 6749 5031 6783
rect 5031 6749 5040 6783
rect 4988 6740 5040 6749
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 3424 6604 3476 6656
rect 4620 6647 4672 6656
rect 4620 6613 4629 6647
rect 4629 6613 4663 6647
rect 4663 6613 4672 6647
rect 4620 6604 4672 6613
rect 5540 6672 5592 6724
rect 6000 6672 6052 6724
rect 5448 6604 5500 6656
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 2136 6400 2188 6452
rect 4620 6400 4672 6452
rect 4896 6400 4948 6452
rect 5448 6400 5500 6452
rect 5540 6400 5592 6452
rect 940 6264 992 6316
rect 3240 6332 3292 6384
rect 3424 6332 3476 6384
rect 4712 6332 4764 6384
rect 5356 6375 5408 6384
rect 5356 6341 5365 6375
rect 5365 6341 5399 6375
rect 5399 6341 5408 6375
rect 5356 6332 5408 6341
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 2780 6264 2832 6273
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 2596 6196 2648 6248
rect 3884 6196 3936 6248
rect 4528 6196 4580 6248
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 2228 6103 2280 6112
rect 2228 6069 2237 6103
rect 2237 6069 2271 6103
rect 2271 6069 2280 6103
rect 2228 6060 2280 6069
rect 3056 6060 3108 6112
rect 5908 6307 5960 6316
rect 5908 6273 5917 6307
rect 5917 6273 5951 6307
rect 5951 6273 5960 6307
rect 5908 6264 5960 6273
rect 6000 6128 6052 6180
rect 3792 6060 3844 6112
rect 3976 6060 4028 6112
rect 5356 6060 5408 6112
rect 2350 5958 2402 6010
rect 2414 5958 2466 6010
rect 2478 5958 2530 6010
rect 2542 5958 2594 6010
rect 2606 5958 2658 6010
rect 1860 5856 1912 5908
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 3792 5899 3844 5908
rect 3792 5865 3801 5899
rect 3801 5865 3835 5899
rect 3835 5865 3844 5899
rect 3792 5856 3844 5865
rect 4436 5856 4488 5908
rect 4528 5856 4580 5908
rect 4620 5856 4672 5908
rect 2228 5720 2280 5772
rect 3056 5720 3108 5772
rect 3516 5720 3568 5772
rect 3976 5720 4028 5772
rect 3884 5652 3936 5704
rect 4344 5652 4396 5704
rect 4988 5788 5040 5840
rect 5540 5788 5592 5840
rect 4896 5695 4948 5704
rect 4896 5661 4905 5695
rect 4905 5661 4939 5695
rect 4939 5661 4948 5695
rect 4896 5652 4948 5661
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 5448 5652 5500 5704
rect 2964 5584 3016 5636
rect 4160 5627 4212 5636
rect 4160 5593 4169 5627
rect 4169 5593 4203 5627
rect 4203 5593 4212 5627
rect 4160 5584 4212 5593
rect 4068 5516 4120 5568
rect 4712 5516 4764 5568
rect 4804 5516 4856 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 4344 5312 4396 5364
rect 4620 5312 4672 5364
rect 4804 5312 4856 5364
rect 5080 5312 5132 5364
rect 2872 5244 2924 5296
rect 4160 5244 4212 5296
rect 4344 5219 4396 5228
rect 4344 5185 4353 5219
rect 4353 5185 4387 5219
rect 4387 5185 4396 5219
rect 4344 5176 4396 5185
rect 4620 5176 4672 5228
rect 4712 5108 4764 5160
rect 5356 5176 5408 5228
rect 6644 5176 6696 5228
rect 5264 5108 5316 5160
rect 7012 5108 7064 5160
rect 5080 5040 5132 5092
rect 5172 5040 5224 5092
rect 940 4972 992 5024
rect 6828 4972 6880 5024
rect 2350 4870 2402 4922
rect 2414 4870 2466 4922
rect 2478 4870 2530 4922
rect 2542 4870 2594 4922
rect 2606 4870 2658 4922
rect 1032 4768 1084 4820
rect 4988 4768 5040 4820
rect 6920 4768 6972 4820
rect 2228 4675 2280 4684
rect 2228 4641 2237 4675
rect 2237 4641 2271 4675
rect 2271 4641 2280 4675
rect 2228 4632 2280 4641
rect 3332 4632 3384 4684
rect 5540 4675 5592 4684
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 2136 4564 2188 4616
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 2780 4564 2832 4616
rect 3608 4496 3660 4548
rect 4896 4496 4948 4548
rect 5172 4564 5224 4616
rect 5816 4496 5868 4548
rect 6000 4496 6052 4548
rect 4160 4428 4212 4480
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 4160 4224 4212 4276
rect 5264 4224 5316 4276
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 2688 4156 2740 4208
rect 2780 4088 2832 4140
rect 3792 4131 3844 4140
rect 3792 4097 3801 4131
rect 3801 4097 3835 4131
rect 3835 4097 3844 4131
rect 3792 4088 3844 4097
rect 3884 4131 3936 4140
rect 3884 4097 3893 4131
rect 3893 4097 3927 4131
rect 3927 4097 3936 4131
rect 3884 4088 3936 4097
rect 3976 4088 4028 4140
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 1952 4063 2004 4072
rect 1952 4029 1961 4063
rect 1961 4029 1995 4063
rect 1995 4029 2004 4063
rect 1952 4020 2004 4029
rect 3516 4020 3568 4072
rect 4068 4020 4120 4072
rect 2780 3952 2832 4004
rect 2228 3884 2280 3936
rect 2504 3884 2556 3936
rect 4344 3952 4396 4004
rect 2964 3884 3016 3936
rect 3056 3927 3108 3936
rect 3056 3893 3065 3927
rect 3065 3893 3099 3927
rect 3099 3893 3108 3927
rect 3056 3884 3108 3893
rect 3240 3927 3292 3936
rect 3240 3893 3249 3927
rect 3249 3893 3283 3927
rect 3283 3893 3292 3927
rect 3240 3884 3292 3893
rect 4068 3927 4120 3936
rect 4068 3893 4077 3927
rect 4077 3893 4111 3927
rect 4111 3893 4120 3927
rect 4068 3884 4120 3893
rect 4620 3995 4672 4004
rect 4620 3961 4629 3995
rect 4629 3961 4663 3995
rect 4663 3961 4672 3995
rect 4620 3952 4672 3961
rect 5908 4088 5960 4140
rect 6644 4088 6696 4140
rect 5724 4063 5776 4072
rect 5724 4029 5733 4063
rect 5733 4029 5767 4063
rect 5767 4029 5776 4063
rect 5724 4020 5776 4029
rect 5632 3952 5684 4004
rect 6828 4020 6880 4072
rect 5264 3884 5316 3936
rect 5448 3884 5500 3936
rect 2350 3782 2402 3834
rect 2414 3782 2466 3834
rect 2478 3782 2530 3834
rect 2542 3782 2594 3834
rect 2606 3782 2658 3834
rect 1860 3680 1912 3732
rect 2228 3680 2280 3732
rect 2596 3612 2648 3664
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 4068 3680 4120 3732
rect 2780 3612 2832 3664
rect 3056 3612 3108 3664
rect 3240 3612 3292 3664
rect 3976 3612 4028 3664
rect 4804 3680 4856 3732
rect 5080 3680 5132 3732
rect 5540 3723 5592 3732
rect 5540 3689 5549 3723
rect 5549 3689 5583 3723
rect 5583 3689 5592 3723
rect 5540 3680 5592 3689
rect 5632 3680 5684 3732
rect 5724 3680 5776 3732
rect 940 3476 992 3528
rect 2320 3587 2372 3596
rect 2320 3553 2329 3587
rect 2329 3553 2363 3587
rect 2363 3553 2372 3587
rect 2320 3544 2372 3553
rect 2044 3476 2096 3528
rect 2504 3408 2556 3460
rect 2872 3476 2924 3528
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 3240 3476 3292 3528
rect 4528 3544 4580 3596
rect 5264 3544 5316 3596
rect 7012 3587 7064 3596
rect 7012 3553 7021 3587
rect 7021 3553 7055 3587
rect 7055 3553 7064 3587
rect 7012 3544 7064 3553
rect 3608 3408 3660 3460
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 4252 3476 4304 3528
rect 2228 3340 2280 3392
rect 2964 3383 3016 3392
rect 2964 3349 2973 3383
rect 2973 3349 3007 3383
rect 3007 3349 3016 3383
rect 2964 3340 3016 3349
rect 3056 3340 3108 3392
rect 4988 3519 5040 3528
rect 4988 3485 4997 3519
rect 4997 3485 5031 3519
rect 5031 3485 5040 3519
rect 4988 3476 5040 3485
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 5448 3519 5500 3528
rect 5448 3485 5457 3519
rect 5457 3485 5491 3519
rect 5491 3485 5500 3519
rect 5448 3476 5500 3485
rect 5540 3476 5592 3528
rect 6552 3476 6604 3528
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 2228 3136 2280 3188
rect 2872 3136 2924 3188
rect 3424 3136 3476 3188
rect 3792 3179 3844 3188
rect 3792 3145 3801 3179
rect 3801 3145 3835 3179
rect 3835 3145 3844 3179
rect 3792 3136 3844 3145
rect 4068 3136 4120 3188
rect 4528 3136 4580 3188
rect 940 3000 992 3052
rect 4988 3136 5040 3188
rect 5172 3136 5224 3188
rect 6920 3136 6972 3188
rect 2688 2864 2740 2916
rect 3516 2864 3568 2916
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 4896 3043 4948 3052
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 2136 2796 2188 2848
rect 2504 2796 2556 2848
rect 6552 2839 6604 2848
rect 6552 2805 6561 2839
rect 6561 2805 6595 2839
rect 6595 2805 6604 2839
rect 6552 2796 6604 2805
rect 2350 2694 2402 2746
rect 2414 2694 2466 2746
rect 2478 2694 2530 2746
rect 2542 2694 2594 2746
rect 2606 2694 2658 2746
rect 5816 2592 5868 2644
rect 6644 2456 6696 2508
rect 6552 2388 6604 2440
rect 6828 2431 6880 2440
rect 6828 2397 6837 2431
rect 6837 2397 6871 2431
rect 6871 2397 6880 2431
rect 6828 2388 6880 2397
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
<< metal2 >>
rect 5170 9832 5226 10632
rect 2350 8188 2658 8197
rect 2350 8186 2356 8188
rect 2412 8186 2436 8188
rect 2492 8186 2516 8188
rect 2572 8186 2596 8188
rect 2652 8186 2658 8188
rect 2412 8134 2414 8186
rect 2594 8134 2596 8186
rect 2350 8132 2356 8134
rect 2412 8132 2436 8134
rect 2492 8132 2516 8134
rect 2572 8132 2596 8134
rect 2652 8132 2658 8134
rect 2350 8123 2658 8132
rect 5184 7886 5212 9832
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 1492 7812 1544 7818
rect 1492 7754 1544 7760
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 1306 7576 1362 7585
rect 1306 7511 1308 7520
rect 1360 7511 1362 7520
rect 1308 7482 1360 7488
rect 1504 6905 1532 7754
rect 2148 7478 2176 7754
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 1872 6662 1900 7142
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 940 6316 992 6322
rect 940 6258 992 6264
rect 952 6225 980 6258
rect 938 6216 994 6225
rect 938 6151 994 6160
rect 1872 5914 1900 6598
rect 1964 6118 1992 7414
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2350 7100 2658 7109
rect 2350 7098 2356 7100
rect 2412 7098 2436 7100
rect 2492 7098 2516 7100
rect 2572 7098 2596 7100
rect 2652 7098 2658 7100
rect 2412 7046 2414 7098
rect 2594 7046 2596 7098
rect 2350 7044 2356 7046
rect 2412 7044 2436 7046
rect 2492 7044 2516 7046
rect 2572 7044 2596 7046
rect 2652 7044 2658 7046
rect 2350 7035 2658 7044
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1030 5536 1086 5545
rect 1030 5471 1086 5480
rect 940 5024 992 5030
rect 940 4966 992 4972
rect 952 4865 980 4966
rect 938 4856 994 4865
rect 1044 4826 1072 5471
rect 938 4791 994 4800
rect 1032 4820 1084 4826
rect 1032 4762 1084 4768
rect 1398 4176 1454 4185
rect 1398 4111 1400 4120
rect 1452 4111 1454 4120
rect 1860 4140 1912 4146
rect 1400 4082 1452 4088
rect 1860 4082 1912 4088
rect 1872 3738 1900 4082
rect 1964 4078 1992 6054
rect 2148 4622 2176 6394
rect 2516 6322 2544 6938
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2608 6254 2636 6666
rect 2792 6322 2820 7142
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 3436 6390 3464 6598
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3424 6384 3476 6390
rect 3424 6326 3476 6332
rect 2780 6316 2832 6322
rect 2964 6316 3016 6322
rect 2832 6276 2912 6304
rect 2780 6258 2832 6264
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2240 5778 2268 6054
rect 2350 6012 2658 6021
rect 2350 6010 2356 6012
rect 2412 6010 2436 6012
rect 2492 6010 2516 6012
rect 2572 6010 2596 6012
rect 2652 6010 2658 6012
rect 2412 5958 2414 6010
rect 2594 5958 2596 6010
rect 2350 5956 2356 5958
rect 2412 5956 2436 5958
rect 2492 5956 2516 5958
rect 2572 5956 2596 5958
rect 2652 5956 2658 5958
rect 2350 5947 2658 5956
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 2240 4690 2268 5714
rect 2884 5302 2912 6276
rect 2964 6258 3016 6264
rect 2976 5642 3004 6258
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3068 5778 3096 6054
rect 3252 5914 3280 6326
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2350 4924 2658 4933
rect 2350 4922 2356 4924
rect 2412 4922 2436 4924
rect 2492 4922 2516 4924
rect 2572 4922 2596 4924
rect 2652 4922 2658 4924
rect 2412 4870 2414 4922
rect 2594 4870 2596 4922
rect 2350 4868 2356 4870
rect 2412 4868 2436 4870
rect 2492 4868 2516 4870
rect 2572 4868 2596 4870
rect 2652 4868 2658 4870
rect 2350 4859 2658 4868
rect 2884 4706 2912 5238
rect 3436 4706 3464 6326
rect 3896 6254 3924 7754
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4172 6798 4200 6938
rect 5276 6866 5304 7142
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3804 5914 3832 6054
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 2700 4678 2912 4706
rect 3344 4690 3464 4706
rect 3332 4684 3464 4690
rect 2136 4616 2188 4622
rect 2056 4576 2136 4604
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2056 3534 2084 4576
rect 2136 4558 2188 4564
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2332 4026 2360 4558
rect 2700 4214 2728 4678
rect 3384 4678 3464 4684
rect 3332 4626 3384 4632
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2688 4208 2740 4214
rect 2688 4150 2740 4156
rect 2148 3998 2452 4026
rect 940 3528 992 3534
rect 938 3496 940 3505
rect 2044 3528 2096 3534
rect 992 3496 994 3505
rect 2044 3470 2096 3476
rect 938 3431 994 3440
rect 940 3052 992 3058
rect 940 2994 992 3000
rect 952 2825 980 2994
rect 2148 2854 2176 3998
rect 2228 3936 2280 3942
rect 2424 3924 2452 3998
rect 2504 3936 2556 3942
rect 2424 3896 2504 3924
rect 2228 3878 2280 3884
rect 2504 3878 2556 3884
rect 2240 3738 2268 3878
rect 2350 3836 2658 3845
rect 2350 3834 2356 3836
rect 2412 3834 2436 3836
rect 2492 3834 2516 3836
rect 2572 3834 2596 3836
rect 2652 3834 2658 3836
rect 2412 3782 2414 3834
rect 2594 3782 2596 3834
rect 2350 3780 2356 3782
rect 2412 3780 2436 3782
rect 2492 3780 2516 3782
rect 2572 3780 2596 3782
rect 2652 3780 2658 3782
rect 2350 3771 2658 3780
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2596 3664 2648 3670
rect 2318 3632 2374 3641
rect 2596 3606 2648 3612
rect 2318 3567 2320 3576
rect 2372 3567 2374 3576
rect 2320 3538 2372 3544
rect 2608 3505 2636 3606
rect 2594 3496 2650 3505
rect 2504 3460 2556 3466
rect 2594 3431 2650 3440
rect 2504 3402 2556 3408
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2240 3194 2268 3334
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2516 2854 2544 3402
rect 2700 2922 2728 4150
rect 2792 4146 2820 4558
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2792 4010 2820 4082
rect 3528 4078 3556 5714
rect 3896 5710 3924 6190
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5778 4016 6054
rect 4066 5944 4122 5953
rect 4448 5914 4476 6734
rect 4540 6254 4568 6734
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4632 6458 4660 6598
rect 4620 6452 4672 6458
rect 4896 6452 4948 6458
rect 4620 6394 4672 6400
rect 4816 6412 4896 6440
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4540 5914 4568 6190
rect 4618 5944 4674 5953
rect 4066 5879 4122 5888
rect 4436 5908 4488 5914
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 4080 5574 4108 5879
rect 4436 5850 4488 5856
rect 4528 5908 4580 5914
rect 4618 5879 4620 5888
rect 4528 5850 4580 5856
rect 4672 5879 4674 5888
rect 4620 5850 4672 5856
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4172 5302 4200 5578
rect 4356 5370 4384 5646
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 3608 4548 3660 4554
rect 3608 4490 3660 4496
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2792 3670 2820 3946
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2884 3194 2912 3470
rect 2976 3398 3004 3878
rect 3068 3670 3096 3878
rect 3252 3670 3280 3878
rect 3056 3664 3108 3670
rect 3240 3664 3292 3670
rect 3056 3606 3108 3612
rect 3238 3632 3240 3641
rect 3292 3632 3294 3641
rect 3238 3567 3294 3576
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 3240 3528 3292 3534
rect 3292 3488 3464 3516
rect 3240 3470 3292 3476
rect 3068 3398 3096 3470
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 3436 3194 3464 3488
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3528 2922 3556 4014
rect 3620 3466 3648 4490
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4172 4282 4200 4422
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 3608 3460 3660 3466
rect 3608 3402 3660 3408
rect 3804 3194 3832 4082
rect 3896 3738 3924 4082
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3988 3670 4016 4082
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4080 3942 4108 4014
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3738 4108 3878
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3988 3505 4016 3606
rect 4264 3534 4292 4082
rect 4356 4010 4384 5170
rect 4448 5114 4476 5850
rect 4724 5760 4752 6326
rect 4632 5732 4752 5760
rect 4632 5370 4660 5732
rect 4816 5658 4844 6412
rect 4896 6394 4948 6400
rect 5000 5846 5028 6734
rect 4988 5840 5040 5846
rect 4988 5782 5040 5788
rect 4724 5630 4844 5658
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4724 5574 4752 5630
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4632 5234 4660 5306
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4724 5166 4752 5510
rect 4816 5370 4844 5510
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4712 5160 4764 5166
rect 4448 5086 4660 5114
rect 4764 5120 4844 5148
rect 4712 5102 4764 5108
rect 4632 4010 4660 5086
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4816 3890 4844 5120
rect 4908 4554 4936 5646
rect 5000 4826 5028 5782
rect 5276 5710 5304 6802
rect 5368 6390 5396 6802
rect 5460 6662 5488 7686
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6840 6905 6868 7142
rect 6826 6896 6882 6905
rect 6826 6831 6882 6840
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 6000 6724 6052 6730
rect 6000 6666 6052 6672
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5460 6458 5488 6598
rect 5552 6458 5580 6666
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5092 5098 5120 5306
rect 5368 5234 5396 6054
rect 5460 5710 5488 6394
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 4816 3862 4936 3890
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4068 3528 4120 3534
rect 3974 3496 4030 3505
rect 4068 3470 4120 3476
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 3974 3431 4030 3440
rect 4080 3194 4108 3470
rect 4540 3194 4568 3538
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4816 3058 4844 3674
rect 4908 3058 4936 3862
rect 5092 3738 5120 5034
rect 5184 4622 5212 5034
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5276 4282 5304 5102
rect 5552 4690 5580 5782
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5276 3602 5304 3878
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5460 3534 5488 3878
rect 5644 3738 5672 3946
rect 5736 3738 5764 4014
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5552 3534 5580 3674
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5000 3194 5028 3470
rect 5184 3194 5212 3470
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 2136 2848 2188 2854
rect 938 2816 994 2825
rect 2136 2790 2188 2796
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 938 2751 994 2760
rect 2350 2748 2658 2757
rect 2350 2746 2356 2748
rect 2412 2746 2436 2748
rect 2492 2746 2516 2748
rect 2572 2746 2596 2748
rect 2652 2746 2658 2748
rect 2412 2694 2414 2746
rect 2594 2694 2596 2746
rect 2350 2692 2356 2694
rect 2412 2692 2436 2694
rect 2492 2692 2516 2694
rect 2572 2692 2596 2694
rect 2652 2692 2658 2694
rect 2350 2683 2658 2692
rect 5828 2650 5856 4490
rect 5920 4146 5948 6258
rect 6012 6186 6040 6666
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 6012 4554 6040 6122
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 6656 4146 6684 5170
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6564 2854 6592 3470
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 6564 2446 6592 2790
rect 6656 2514 6684 4082
rect 6840 4078 6868 4966
rect 6932 4826 6960 7346
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7024 4865 7052 5102
rect 7010 4856 7066 4865
rect 6920 4820 6972 4826
rect 7010 4791 7066 4800
rect 6920 4762 6972 4768
rect 7010 4176 7066 4185
rect 7010 4111 7066 4120
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 6840 2446 6868 4014
rect 7024 3602 7052 4111
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6918 3496 6974 3505
rect 6918 3431 6974 3440
rect 6932 3194 6960 3431
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
<< via2 >>
rect 2356 8186 2412 8188
rect 2436 8186 2492 8188
rect 2516 8186 2572 8188
rect 2596 8186 2652 8188
rect 2356 8134 2402 8186
rect 2402 8134 2412 8186
rect 2436 8134 2466 8186
rect 2466 8134 2478 8186
rect 2478 8134 2492 8186
rect 2516 8134 2530 8186
rect 2530 8134 2542 8186
rect 2542 8134 2572 8186
rect 2596 8134 2606 8186
rect 2606 8134 2652 8186
rect 2356 8132 2412 8134
rect 2436 8132 2492 8134
rect 2516 8132 2572 8134
rect 2596 8132 2652 8134
rect 1306 7540 1362 7576
rect 1306 7520 1308 7540
rect 1308 7520 1360 7540
rect 1360 7520 1362 7540
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 1490 6840 1546 6896
rect 938 6160 994 6216
rect 2356 7098 2412 7100
rect 2436 7098 2492 7100
rect 2516 7098 2572 7100
rect 2596 7098 2652 7100
rect 2356 7046 2402 7098
rect 2402 7046 2412 7098
rect 2436 7046 2466 7098
rect 2466 7046 2478 7098
rect 2478 7046 2492 7098
rect 2516 7046 2530 7098
rect 2530 7046 2542 7098
rect 2542 7046 2572 7098
rect 2596 7046 2606 7098
rect 2606 7046 2652 7098
rect 2356 7044 2412 7046
rect 2436 7044 2492 7046
rect 2516 7044 2572 7046
rect 2596 7044 2652 7046
rect 1030 5480 1086 5536
rect 938 4800 994 4856
rect 1398 4140 1454 4176
rect 1398 4120 1400 4140
rect 1400 4120 1452 4140
rect 1452 4120 1454 4140
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 2356 6010 2412 6012
rect 2436 6010 2492 6012
rect 2516 6010 2572 6012
rect 2596 6010 2652 6012
rect 2356 5958 2402 6010
rect 2402 5958 2412 6010
rect 2436 5958 2466 6010
rect 2466 5958 2478 6010
rect 2478 5958 2492 6010
rect 2516 5958 2530 6010
rect 2530 5958 2542 6010
rect 2542 5958 2572 6010
rect 2596 5958 2606 6010
rect 2606 5958 2652 6010
rect 2356 5956 2412 5958
rect 2436 5956 2492 5958
rect 2516 5956 2572 5958
rect 2596 5956 2652 5958
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 2356 4922 2412 4924
rect 2436 4922 2492 4924
rect 2516 4922 2572 4924
rect 2596 4922 2652 4924
rect 2356 4870 2402 4922
rect 2402 4870 2412 4922
rect 2436 4870 2466 4922
rect 2466 4870 2478 4922
rect 2478 4870 2492 4922
rect 2516 4870 2530 4922
rect 2530 4870 2542 4922
rect 2542 4870 2572 4922
rect 2596 4870 2606 4922
rect 2606 4870 2652 4922
rect 2356 4868 2412 4870
rect 2436 4868 2492 4870
rect 2516 4868 2572 4870
rect 2596 4868 2652 4870
rect 938 3476 940 3496
rect 940 3476 992 3496
rect 992 3476 994 3496
rect 938 3440 994 3476
rect 2356 3834 2412 3836
rect 2436 3834 2492 3836
rect 2516 3834 2572 3836
rect 2596 3834 2652 3836
rect 2356 3782 2402 3834
rect 2402 3782 2412 3834
rect 2436 3782 2466 3834
rect 2466 3782 2478 3834
rect 2478 3782 2492 3834
rect 2516 3782 2530 3834
rect 2530 3782 2542 3834
rect 2542 3782 2572 3834
rect 2596 3782 2606 3834
rect 2606 3782 2652 3834
rect 2356 3780 2412 3782
rect 2436 3780 2492 3782
rect 2516 3780 2572 3782
rect 2596 3780 2652 3782
rect 2318 3596 2374 3632
rect 2318 3576 2320 3596
rect 2320 3576 2372 3596
rect 2372 3576 2374 3596
rect 2594 3440 2650 3496
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 4066 5888 4122 5944
rect 4618 5908 4674 5944
rect 4618 5888 4620 5908
rect 4620 5888 4672 5908
rect 4672 5888 4674 5908
rect 3238 3612 3240 3632
rect 3240 3612 3292 3632
rect 3292 3612 3294 3632
rect 3238 3576 3294 3612
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 6826 6840 6882 6896
rect 3974 3440 4030 3496
rect 938 2760 994 2816
rect 2356 2746 2412 2748
rect 2436 2746 2492 2748
rect 2516 2746 2572 2748
rect 2596 2746 2652 2748
rect 2356 2694 2402 2746
rect 2402 2694 2412 2746
rect 2436 2694 2466 2746
rect 2466 2694 2478 2746
rect 2478 2694 2492 2746
rect 2516 2694 2530 2746
rect 2530 2694 2542 2746
rect 2542 2694 2572 2746
rect 2596 2694 2606 2746
rect 2606 2694 2652 2746
rect 2356 2692 2412 2694
rect 2436 2692 2492 2694
rect 2516 2692 2572 2694
rect 2596 2692 2652 2694
rect 7010 4800 7066 4856
rect 7010 4120 7066 4176
rect 6918 3440 6974 3496
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
<< metal3 >>
rect 2346 8192 2662 8193
rect 2346 8128 2352 8192
rect 2416 8128 2432 8192
rect 2496 8128 2512 8192
rect 2576 8128 2592 8192
rect 2656 8128 2662 8192
rect 2346 8127 2662 8128
rect 3006 7648 3322 7649
rect 0 7578 800 7608
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 1301 7578 1367 7581
rect 0 7576 1367 7578
rect 0 7520 1306 7576
rect 1362 7520 1367 7576
rect 0 7518 1367 7520
rect 0 7488 800 7518
rect 1301 7515 1367 7518
rect 2346 7104 2662 7105
rect 2346 7040 2352 7104
rect 2416 7040 2432 7104
rect 2496 7040 2512 7104
rect 2576 7040 2592 7104
rect 2656 7040 2662 7104
rect 2346 7039 2662 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 6821 6898 6887 6901
rect 7688 6898 8488 6928
rect 6821 6896 8488 6898
rect 6821 6840 6826 6896
rect 6882 6840 8488 6896
rect 6821 6838 8488 6840
rect 6821 6835 6887 6838
rect 7688 6808 8488 6838
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 0 6218 800 6248
rect 933 6218 999 6221
rect 0 6216 999 6218
rect 0 6160 938 6216
rect 994 6160 999 6216
rect 0 6158 999 6160
rect 0 6128 800 6158
rect 933 6155 999 6158
rect 2346 6016 2662 6017
rect 2346 5952 2352 6016
rect 2416 5952 2432 6016
rect 2496 5952 2512 6016
rect 2576 5952 2592 6016
rect 2656 5952 2662 6016
rect 2346 5951 2662 5952
rect 4061 5946 4127 5949
rect 4613 5946 4679 5949
rect 4061 5944 4679 5946
rect 4061 5888 4066 5944
rect 4122 5888 4618 5944
rect 4674 5888 4679 5944
rect 4061 5886 4679 5888
rect 4061 5883 4127 5886
rect 4613 5883 4679 5886
rect 0 5538 800 5568
rect 1025 5538 1091 5541
rect 0 5536 1091 5538
rect 0 5480 1030 5536
rect 1086 5480 1091 5536
rect 0 5478 1091 5480
rect 0 5448 800 5478
rect 1025 5475 1091 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 2346 4928 2662 4929
rect 0 4858 800 4888
rect 2346 4864 2352 4928
rect 2416 4864 2432 4928
rect 2496 4864 2512 4928
rect 2576 4864 2592 4928
rect 2656 4864 2662 4928
rect 2346 4863 2662 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 7005 4858 7071 4861
rect 7688 4858 8488 4888
rect 7005 4856 8488 4858
rect 7005 4800 7010 4856
rect 7066 4800 8488 4856
rect 7005 4798 8488 4800
rect 7005 4795 7071 4798
rect 7688 4768 8488 4798
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 0 4178 800 4208
rect 1393 4178 1459 4181
rect 0 4176 1459 4178
rect 0 4120 1398 4176
rect 1454 4120 1459 4176
rect 0 4118 1459 4120
rect 0 4088 800 4118
rect 1393 4115 1459 4118
rect 7005 4178 7071 4181
rect 7688 4178 8488 4208
rect 7005 4176 8488 4178
rect 7005 4120 7010 4176
rect 7066 4120 8488 4176
rect 7005 4118 8488 4120
rect 7005 4115 7071 4118
rect 7688 4088 8488 4118
rect 2346 3840 2662 3841
rect 2346 3776 2352 3840
rect 2416 3776 2432 3840
rect 2496 3776 2512 3840
rect 2576 3776 2592 3840
rect 2656 3776 2662 3840
rect 2346 3775 2662 3776
rect 2313 3634 2379 3637
rect 3233 3634 3299 3637
rect 2313 3632 3299 3634
rect 2313 3576 2318 3632
rect 2374 3576 3238 3632
rect 3294 3576 3299 3632
rect 2313 3574 3299 3576
rect 2313 3571 2379 3574
rect 3233 3571 3299 3574
rect 0 3498 800 3528
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 2589 3498 2655 3501
rect 3969 3498 4035 3501
rect 2589 3496 4035 3498
rect 2589 3440 2594 3496
rect 2650 3440 3974 3496
rect 4030 3440 4035 3496
rect 2589 3438 4035 3440
rect 2589 3435 2655 3438
rect 3969 3435 4035 3438
rect 6913 3498 6979 3501
rect 7688 3498 8488 3528
rect 6913 3496 8488 3498
rect 6913 3440 6918 3496
rect 6974 3440 8488 3496
rect 6913 3438 8488 3440
rect 6913 3435 6979 3438
rect 7688 3408 8488 3438
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 2346 2752 2662 2753
rect 2346 2688 2352 2752
rect 2416 2688 2432 2752
rect 2496 2688 2512 2752
rect 2576 2688 2592 2752
rect 2656 2688 2662 2752
rect 2346 2687 2662 2688
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
<< via3 >>
rect 2352 8188 2416 8192
rect 2352 8132 2356 8188
rect 2356 8132 2412 8188
rect 2412 8132 2416 8188
rect 2352 8128 2416 8132
rect 2432 8188 2496 8192
rect 2432 8132 2436 8188
rect 2436 8132 2492 8188
rect 2492 8132 2496 8188
rect 2432 8128 2496 8132
rect 2512 8188 2576 8192
rect 2512 8132 2516 8188
rect 2516 8132 2572 8188
rect 2572 8132 2576 8188
rect 2512 8128 2576 8132
rect 2592 8188 2656 8192
rect 2592 8132 2596 8188
rect 2596 8132 2652 8188
rect 2652 8132 2656 8188
rect 2592 8128 2656 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 2352 7100 2416 7104
rect 2352 7044 2356 7100
rect 2356 7044 2412 7100
rect 2412 7044 2416 7100
rect 2352 7040 2416 7044
rect 2432 7100 2496 7104
rect 2432 7044 2436 7100
rect 2436 7044 2492 7100
rect 2492 7044 2496 7100
rect 2432 7040 2496 7044
rect 2512 7100 2576 7104
rect 2512 7044 2516 7100
rect 2516 7044 2572 7100
rect 2572 7044 2576 7100
rect 2512 7040 2576 7044
rect 2592 7100 2656 7104
rect 2592 7044 2596 7100
rect 2596 7044 2652 7100
rect 2652 7044 2656 7100
rect 2592 7040 2656 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 2352 6012 2416 6016
rect 2352 5956 2356 6012
rect 2356 5956 2412 6012
rect 2412 5956 2416 6012
rect 2352 5952 2416 5956
rect 2432 6012 2496 6016
rect 2432 5956 2436 6012
rect 2436 5956 2492 6012
rect 2492 5956 2496 6012
rect 2432 5952 2496 5956
rect 2512 6012 2576 6016
rect 2512 5956 2516 6012
rect 2516 5956 2572 6012
rect 2572 5956 2576 6012
rect 2512 5952 2576 5956
rect 2592 6012 2656 6016
rect 2592 5956 2596 6012
rect 2596 5956 2652 6012
rect 2652 5956 2656 6012
rect 2592 5952 2656 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 2352 4924 2416 4928
rect 2352 4868 2356 4924
rect 2356 4868 2412 4924
rect 2412 4868 2416 4924
rect 2352 4864 2416 4868
rect 2432 4924 2496 4928
rect 2432 4868 2436 4924
rect 2436 4868 2492 4924
rect 2492 4868 2496 4924
rect 2432 4864 2496 4868
rect 2512 4924 2576 4928
rect 2512 4868 2516 4924
rect 2516 4868 2572 4924
rect 2572 4868 2576 4924
rect 2512 4864 2576 4868
rect 2592 4924 2656 4928
rect 2592 4868 2596 4924
rect 2596 4868 2652 4924
rect 2652 4868 2656 4924
rect 2592 4864 2656 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 2352 3836 2416 3840
rect 2352 3780 2356 3836
rect 2356 3780 2412 3836
rect 2412 3780 2416 3836
rect 2352 3776 2416 3780
rect 2432 3836 2496 3840
rect 2432 3780 2436 3836
rect 2436 3780 2492 3836
rect 2492 3780 2496 3836
rect 2432 3776 2496 3780
rect 2512 3836 2576 3840
rect 2512 3780 2516 3836
rect 2516 3780 2572 3836
rect 2572 3780 2576 3836
rect 2512 3776 2576 3780
rect 2592 3836 2656 3840
rect 2592 3780 2596 3836
rect 2596 3780 2652 3836
rect 2652 3780 2656 3836
rect 2592 3776 2656 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 2352 2748 2416 2752
rect 2352 2692 2356 2748
rect 2356 2692 2412 2748
rect 2412 2692 2416 2748
rect 2352 2688 2416 2692
rect 2432 2748 2496 2752
rect 2432 2692 2436 2748
rect 2436 2692 2492 2748
rect 2492 2692 2496 2748
rect 2432 2688 2496 2692
rect 2512 2748 2576 2752
rect 2512 2692 2516 2748
rect 2516 2692 2572 2748
rect 2572 2692 2576 2748
rect 2512 2688 2576 2692
rect 2592 2748 2656 2752
rect 2592 2692 2596 2748
rect 2596 2692 2652 2748
rect 2652 2692 2656 2748
rect 2592 2688 2656 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
<< metal4 >>
rect 2344 8192 2664 8208
rect 2344 8128 2352 8192
rect 2416 8128 2432 8192
rect 2496 8128 2512 8192
rect 2576 8128 2592 8192
rect 2656 8128 2664 8192
rect 2344 7104 2664 8128
rect 2344 7040 2352 7104
rect 2416 7040 2432 7104
rect 2496 7040 2512 7104
rect 2576 7040 2592 7104
rect 2656 7040 2664 7104
rect 2344 6016 2664 7040
rect 2344 5952 2352 6016
rect 2416 5952 2432 6016
rect 2496 5952 2512 6016
rect 2576 5952 2592 6016
rect 2656 5952 2664 6016
rect 2344 4928 2664 5952
rect 2344 4864 2352 4928
rect 2416 4864 2432 4928
rect 2496 4864 2512 4928
rect 2576 4864 2592 4928
rect 2656 4864 2664 4928
rect 2344 3840 2664 4864
rect 2344 3776 2352 3840
rect 2416 3776 2432 3840
rect 2496 3776 2512 3840
rect 2576 3776 2592 3840
rect 2656 3776 2664 3840
rect 2344 3694 2664 3776
rect 2344 3458 2386 3694
rect 2622 3458 2664 3694
rect 2344 2752 2664 3458
rect 2344 2688 2352 2752
rect 2416 2688 2432 2752
rect 2496 2688 2512 2752
rect 2576 2688 2592 2752
rect 2656 2688 2664 2752
rect 2344 2128 2664 2688
rect 3004 7648 3324 8208
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4354 3092 4384
rect 3156 4354 3172 4384
rect 3236 4354 3252 4384
rect 3316 4320 3324 4384
rect 3004 4118 3046 4320
rect 3282 4118 3324 4320
rect 3004 3296 3324 4118
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 2128 3324 2144
<< via4 >>
rect 2386 3458 2622 3694
rect 3046 4320 3076 4354
rect 3076 4320 3092 4354
rect 3092 4320 3156 4354
rect 3156 4320 3172 4354
rect 3172 4320 3236 4354
rect 3236 4320 3252 4354
rect 3252 4320 3282 4354
rect 3046 4118 3282 4320
<< metal5 >>
rect 1056 4354 7408 4396
rect 1056 4118 3046 4354
rect 3282 4118 7408 4354
rect 1056 4076 7408 4118
rect 1056 3694 7408 3736
rect 1056 3458 2386 3694
rect 2622 3458 7408 3694
rect 1056 3416 7408 3458
use sky130_fd_sc_hd__or3_1  _37_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2576 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _38_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 5888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _39_
timestamp 1694700623
transform 1 0 3128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _40_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2576 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _41_
timestamp 1694700623
transform 1 0 2208 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _42_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 3680 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _43_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2944 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _44_
timestamp 1694700623
transform -1 0 6900 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _45_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _46_
timestamp 1694700623
transform -1 0 2576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _47_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 2576 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a2111oi_1  _48_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _49_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5428 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _50_
timestamp 1694700623
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _51_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3772 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _52_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4140 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _53_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4416 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _54_
timestamp 1694700623
transform 1 0 4048 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _55_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _56_
timestamp 1694700623
transform 1 0 5428 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _57_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 5336 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _58_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6808 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _59_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_2  _60_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4140 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _61_
timestamp 1694700623
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _62_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 5428 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _63_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _64_
timestamp 1694700623
transform -1 0 4232 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _65_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _66_
timestamp 1694700623
transform -1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _67_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _68_
timestamp 1694700623
transform -1 0 3036 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _69_
timestamp 1694700623
transform -1 0 3680 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _70_
timestamp 1694700623
transform -1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _71_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4324 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _72_
timestamp 1694700623
transform -1 0 6808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _73_
timestamp 1694700623
transform 1 0 6624 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _74_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2944 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _75_
timestamp 1694700623
transform 1 0 1656 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _76_
timestamp 1694700623
transform 1 0 2116 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _77_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4508 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _78_
timestamp 1694700623
transform -1 0 5244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _79_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4968 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _80_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _81_ ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3036 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _82_
timestamp 1694700623
transform 1 0 1380 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _83_
timestamp 1694700623
transform 1 0 5244 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3404 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1694700623
transform -1 0 3220 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1694700623
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_3 ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_11
timestamp 1694700623
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_19
timestamp 1694700623
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 1694700623
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_37
timestamp 1694700623
transform 1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_45
timestamp 1694700623
transform 1 0 5244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_57
timestamp 1694700623
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_64
timestamp 1694700623
transform 1 0 6992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_6 ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1656 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_18 ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2760 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_26
timestamp 1694700623
transform 1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_35
timestamp 1694700623
transform 1 0 4324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_46
timestamp 1694700623
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_63
timestamp 1694700623
transform 1 0 6900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_6
timestamp 1694700623
transform 1 0 1656 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_54
timestamp 1694700623
transform 1 0 6072 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_25 ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1694700623
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_62
timestamp 1694700623
transform 1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_9
timestamp 1694700623
transform 1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_18
timestamp 1694700623
transform 1 0 2760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1694700623
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1694700623
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_44
timestamp 1694700623
transform 1 0 5152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 1694700623
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_11
timestamp 1694700623
transform 1 0 2116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_19
timestamp 1694700623
transform 1 0 2852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_27
timestamp 1694700623
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_62
timestamp 1694700623
transform 1 0 6808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1694700623
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1694700623
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_23
timestamp 1694700623
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1694700623
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_41
timestamp 1694700623
transform 1 0 4876 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_23
timestamp 1694700623
transform 1 0 3220 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_45
timestamp 1694700623
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1694700623
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 1694700623
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_7
timestamp 1694700623
transform 1 0 1748 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_15
timestamp 1694700623
transform 1 0 2484 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_23
timestamp 1694700623
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1694700623
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 1694700623
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_37
timestamp 1694700623
transform 1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_48
timestamp 1694700623
transform 1 0 5520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_57
timestamp 1694700623
transform 1 0 6348 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1694700623
transform 1 0 5244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6256 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input3 ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1694700623
transform -1 0 7084 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1694700623
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1694700623
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1694700623
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap13
timestamp 1694700623
transform 1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output8 ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output9 ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 1694700623
transform -1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1694700623
transform -1 0 2116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 1694700623
transform -1 0 7084 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_11
timestamp 1694700623
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_12
timestamp 1694700623
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_13
timestamp 1694700623
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_14
timestamp 1694700623
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_15
timestamp 1694700623
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_16
timestamp 1694700623
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 7360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_17
timestamp 1694700623
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_18
timestamp 1694700623
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_19
timestamp 1694700623
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 7360 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_20
timestamp 1694700623
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_21
timestamp 1694700623
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 7360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_22 ~/.volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_23
timestamp 1694700623
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_24
timestamp 1694700623
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_25
timestamp 1694700623
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_26
timestamp 1694700623
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_27
timestamp 1694700623
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_28
timestamp 1694700623
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 1694700623
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_30
timestamp 1694700623
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_31
timestamp 1694700623
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_32
timestamp 1694700623
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_33
timestamp 1694700623
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_34
timestamp 1694700623
transform 1 0 6256 0 1 7616
box -38 -48 130 592
<< labels >>
flabel metal4 s 3004 2128 3324 8208 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4076 7408 4396 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2344 2128 2664 8208 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3416 7408 3736 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 5170 9832 5226 10632 0 FreeSans 224 90 0 0 clear
port 2 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 clk
port 3 nsew signal input
flabel metal3 s 7688 3408 8488 3528 0 FreeSans 480 0 0 0 count[0]
port 4 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 count[1]
port 5 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 count[2]
port 6 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 count[3]
port 7 nsew signal tristate
flabel metal3 s 7688 4768 8488 4888 0 FreeSans 480 0 0 0 enable
port 8 nsew signal input
flabel metal3 s 7688 6808 8488 6928 0 FreeSans 480 0 0 0 flag
port 9 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 nRST
port 10 nsew signal input
flabel metal3 s 7688 4088 8488 4208 0 FreeSans 480 0 0 0 rollover[0]
port 11 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 rollover[1]
port 12 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 rollover[2]
port 13 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 rollover[3]
port 14 nsew signal input
rlabel metal1 4232 7616 4232 7616 0 VGND
rlabel metal1 4232 8160 4232 8160 0 VPWR
rlabel metal1 5520 3570 5520 3570 0 _00_
rlabel metal1 5474 3162 5474 3162 0 _01_
rlabel metal2 3266 3757 3266 3757 0 _02_
rlabel viali 3174 3501 3174 3501 0 _03_
rlabel metal1 2990 3502 2990 3502 0 _04_
rlabel metal1 4370 3570 4370 3570 0 _05_
rlabel metal1 4186 2992 4186 2992 0 _06_
rlabel metal1 5290 2992 5290 2992 0 _07_
rlabel metal1 5060 3162 5060 3162 0 _08_
rlabel metal1 2116 3570 2116 3570 0 _09_
rlabel metal1 4094 4148 4094 4148 0 _10_
rlabel metal1 5474 3468 5474 3468 0 _11_
rlabel metal1 5888 3706 5888 3706 0 _12_
rlabel metal2 3910 3910 3910 3910 0 _13_
rlabel metal2 3818 3638 3818 3638 0 _14_
rlabel metal1 4140 3706 4140 3706 0 _15_
rlabel metal1 4278 3162 4278 3162 0 _16_
rlabel metal1 5152 3638 5152 3638 0 _17_
rlabel metal1 6808 4046 6808 4046 0 _18_
rlabel metal1 5244 5202 5244 5202 0 _19_
rlabel metal1 6946 2448 6946 2448 0 _20_
rlabel metal1 6164 4114 6164 4114 0 _21_
rlabel metal1 4232 5882 4232 5882 0 _22_
rlabel viali 4646 5675 4646 5675 0 _23_
rlabel metal2 4186 6868 4186 6868 0 _24_
rlabel metal1 4040 5542 4040 5542 0 _25_
rlabel metal1 2438 6222 2438 6222 0 _26_
rlabel viali 4278 6764 4278 6764 0 _27_
rlabel metal1 3204 5610 3204 5610 0 _28_
rlabel metal1 2162 6324 2162 6324 0 _29_
rlabel metal1 4784 5338 4784 5338 0 _30_
rlabel metal1 5152 4590 5152 4590 0 _31_
rlabel metal1 6256 2618 6256 2618 0 _32_
rlabel metal1 4830 4692 4830 4692 0 _33_
rlabel metal2 4186 4352 4186 4352 0 _34_
rlabel metal1 3450 4692 3450 4692 0 _35_
rlabel metal1 4738 4522 4738 4522 0 _36_
rlabel metal1 5244 7854 5244 7854 0 clear
rlabel metal3 1004 7548 1004 7548 0 clk
rlabel metal1 5106 7174 5106 7174 0 clknet_0_clk
rlabel metal1 1886 6664 1886 6664 0 clknet_1_0__leaf_clk
rlabel metal1 5152 4658 5152 4658 0 clknet_1_1__leaf_clk
rlabel metal1 6532 3162 6532 3162 0 count[0]
rlabel metal3 820 6188 820 6188 0 count[1]
rlabel metal3 866 5508 866 5508 0 count[2]
rlabel metal3 820 4828 820 4828 0 count[3]
rlabel metal1 6624 5134 6624 5134 0 enable
rlabel metal2 6854 7021 6854 7021 0 flag
rlabel metal3 1096 6868 1096 6868 0 nRST
rlabel metal1 5474 6358 5474 6358 0 net1
rlabel metal1 4738 6426 4738 6426 0 net10
rlabel metal1 2530 4148 2530 4148 0 net11
rlabel metal1 6992 4794 6992 4794 0 net12
rlabel metal1 4554 4148 4554 4148 0 net13
rlabel metal1 4784 5202 4784 5202 0 net2
rlabel metal2 2162 7616 2162 7616 0 net3
rlabel metal1 6624 2346 6624 2346 0 net4
rlabel metal1 2622 3468 2622 3468 0 net5
rlabel metal1 2714 3672 2714 3672 0 net6
rlabel metal1 1886 3638 1886 3638 0 net7
rlabel metal2 5382 6596 5382 6596 0 net8
rlabel metal1 2346 6120 2346 6120 0 net9
rlabel metal1 5658 6426 5658 6426 0 next_count\[0\]
rlabel metal2 2254 5372 2254 5372 0 next_count\[1\]
rlabel metal1 3404 6358 3404 6358 0 next_count\[2\]
rlabel metal2 1978 5066 1978 5066 0 next_count\[3\]
rlabel metal2 5566 5236 5566 5236 0 next_flag
rlabel metal2 7038 3859 7038 3859 0 rollover[0]
rlabel metal3 820 2788 820 2788 0 rollover[1]
rlabel metal3 1050 4148 1050 4148 0 rollover[2]
rlabel metal3 820 3468 820 3468 0 rollover[3]
<< properties >>
string FIXED_BBOX 0 0 8488 10632
<< end >>
