VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO flex_counter
  CLASS BLOCK ;
  FOREIGN flex_counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 42.440 BY 53.160 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 15.020 10.640 16.620 41.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 20.380 37.040 21.980 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 11.720 10.640 13.320 41.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 17.080 37.040 18.680 ;
    END
  END VPWR
  PIN clear
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 49.160 26.130 53.160 ;
    END
  END clear
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END clk
  PIN count[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 38.440 17.040 42.440 17.640 ;
    END
  END count[0]
  PIN count[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END count[1]
  PIN count[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END count[2]
  PIN count[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END count[3]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 38.440 23.840 42.440 24.440 ;
    END
  END enable
  PIN flag
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 38.440 34.040 42.440 34.640 ;
    END
  END flag
  PIN nRST
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END nRST
  PIN rollover[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 38.440 20.440 42.440 21.040 ;
    END
  END rollover[0]
  PIN rollover[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END rollover[1]
  PIN rollover[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END rollover[2]
  PIN rollover[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END rollover[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 36.800 40.885 ;
      LAYER met1 ;
        RECT 4.670 10.640 36.800 41.040 ;
      LAYER met2 ;
        RECT 4.690 48.880 25.570 49.160 ;
        RECT 26.410 48.880 35.330 49.160 ;
        RECT 4.690 10.695 35.330 48.880 ;
      LAYER met3 ;
        RECT 4.000 38.440 38.440 40.965 ;
        RECT 4.400 37.040 38.440 38.440 ;
        RECT 4.000 35.040 38.440 37.040 ;
        RECT 4.400 33.640 38.040 35.040 ;
        RECT 4.000 31.640 38.440 33.640 ;
        RECT 4.400 30.240 38.440 31.640 ;
        RECT 4.000 28.240 38.440 30.240 ;
        RECT 4.400 26.840 38.440 28.240 ;
        RECT 4.000 24.840 38.440 26.840 ;
        RECT 4.400 23.440 38.040 24.840 ;
        RECT 4.000 21.440 38.440 23.440 ;
        RECT 4.400 20.040 38.040 21.440 ;
        RECT 4.000 18.040 38.440 20.040 ;
        RECT 4.400 16.640 38.040 18.040 ;
        RECT 4.000 14.640 38.440 16.640 ;
        RECT 4.400 13.240 38.440 14.640 ;
        RECT 4.000 10.715 38.440 13.240 ;
  END
END flex_counter
END LIBRARY

